-- megafunction wizard: %ALTPLL_RECONFIG%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altpll_reconfig 

-- ============================================================
-- File Name: video_pll_reconfig.vhd
-- Megafunction Name(s):
-- 			altpll_reconfig
--
-- Simulation Library Files(s):
-- 			altera_mf;cyclone10lp;lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 22.1std.2 Build 922 07/20/2023 SC Lite Edition
-- ************************************************************


--Copyright (C) 2023  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and any partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details, at
--https://fpgasoftware.intel.com/eula.


--altpll_reconfig CBX_AUTO_BLACKBOX="ALL" device_family="Cyclone 10 LP" init_from_rom="NO" scan_init_file="./Atari800XL/mist/ntsc.mif" busy clock counter_param counter_type data_in data_out pll_areset pll_areset_in pll_configupdate pll_scanclk pll_scanclkena pll_scandata pll_scandataout pll_scandone read_param reconfig reset reset_rom_address rom_address_out rom_data_in write_from_rom write_param write_rom_ena
--VERSION_BEGIN 22.1 cbx_altera_syncram_nd_impl 2023:07:20:14:03:03:SC cbx_altpll_reconfig 2023:07:20:14:03:03:SC cbx_altsyncram 2023:07:20:14:03:03:SC cbx_cycloneii 2023:07:20:14:03:03:SC cbx_lpm_add_sub 2023:07:20:14:03:03:SC cbx_lpm_compare 2023:07:20:14:03:03:SC cbx_lpm_counter 2023:07:20:14:03:03:SC cbx_lpm_decode 2023:07:20:14:03:02:SC cbx_lpm_mux 2023:07:20:14:03:03:SC cbx_mgl 2023:07:20:14:14:26:SC cbx_nadder 2023:07:20:14:03:03:SC cbx_stratix 2023:07:20:14:03:03:SC cbx_stratixii 2023:07:20:14:03:03:SC cbx_stratixiii 2023:07:20:14:03:03:SC cbx_stratixv 2023:07:20:14:03:03:SC cbx_util_mgl 2023:07:20:14:03:03:SC  VERSION_END

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY cyclone10lp;
 USE cyclone10lp.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = altsyncram 1 lpm_add_sub 2 lpm_compare 1 lpm_counter 8 lpm_decode 1 lut 3 reg 102 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  video_pll_reconfig_pllrcfg_2871 IS 
	 PORT 
	 ( 
		 busy	:	OUT  STD_LOGIC;
		 clock	:	IN  STD_LOGIC;
		 counter_param	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0');
		 counter_type	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0');
		 data_in	:	IN  STD_LOGIC_VECTOR (8 DOWNTO 0) := (OTHERS => '0');
		 data_out	:	OUT  STD_LOGIC_VECTOR (8 DOWNTO 0);
		 pll_areset	:	OUT  STD_LOGIC;
		 pll_areset_in	:	IN  STD_LOGIC := '0';
		 pll_configupdate	:	OUT  STD_LOGIC;
		 pll_scanclk	:	OUT  STD_LOGIC;
		 pll_scanclkena	:	OUT  STD_LOGIC;
		 pll_scandata	:	OUT  STD_LOGIC;
		 pll_scandataout	:	IN  STD_LOGIC := '0';
		 pll_scandone	:	IN  STD_LOGIC := '0';
		 read_param	:	IN  STD_LOGIC := '0';
		 reconfig	:	IN  STD_LOGIC := '0';
		 reset	:	IN  STD_LOGIC;
		 reset_rom_address	:	IN  STD_LOGIC := '0';
		 rom_address_out	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 rom_data_in	:	IN  STD_LOGIC := '0';
		 write_from_rom	:	IN  STD_LOGIC := '0';
		 write_param	:	IN  STD_LOGIC := '0';
		 write_rom_ena	:	OUT  STD_LOGIC
	 ); 
 END video_pll_reconfig_pllrcfg_2871;

 ARCHITECTURE RTL OF video_pll_reconfig_pllrcfg_2871 IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "ADV_NETLIST_OPT_ALLOWED=""NEVER_ALLOW"";suppress_da_rule_internal=C106;{-to le_comb10} PLL_SCAN_RECONFIG_COUNTER_REMAP_LCELL=2;{-to le_comb8} PLL_SCAN_RECONFIG_COUNTER_REMAP_LCELL=0;{-to le_comb9} PLL_SCAN_RECONFIG_COUNTER_REMAP_LCELL=1";

	 SIGNAL  wire_altsyncram4_data_a	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altsyncram4_q_a	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_le_comb10_combout	:	STD_LOGIC;
	 SIGNAL  wire_le_comb8_combout	:	STD_LOGIC;
	 SIGNAL  wire_le_comb9_combout	:	STD_LOGIC;
	 SIGNAL	 addr_from_rom	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 addr_from_rom2	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 areset_init_state_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 areset_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 C0_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 C0_ena_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 C1_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 C1_ena_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_C1_ena_state_w_lg_q1786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 C2_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 C2_ena_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_C2_ena_state_w_lg_q1787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 C3_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 C3_ena_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 C4_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 C4_ena_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 configupdate2_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 configupdate3_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_configupdate3_state_w_lg_q1879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 configupdate_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 counter_param_latch_reg	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 counter_type_latch_reg	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 idle_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF idle_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_idle_state_w_lg_w_lg_w_lg_w_lg_q1743w1744w1745w1746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_idle_state_w_lg_w_lg_w_lg_q1743w1744w1745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_idle_state_w_lg_w_lg_q1743w1744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_idle_state_w_lg_q1743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_idle_state_w_lg_q1672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_idle_state_w1747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_idle_state_w_lg_w1747w1748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_idle_state_w_lg_w_lg_w1747w1748w1749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_idle_state_w_lg_w_lg_w_lg_w1747w1748w1749w1750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 nominal_data0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nominal_data1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nominal_data2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nominal_data3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nominal_data4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nominal_data5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nominal_data6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nominal_data7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nominal_data8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nominal_data9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nominal_data10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nominal_data11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nominal_data12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nominal_data13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nominal_data14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nominal_data15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nominal_data16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nominal_data17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_data_nominal_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF read_data_nominal_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_read_data_nominal_state_w_lg_q1772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_data_nominal_state_w_lg_q1686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 read_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF read_data_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_read_data_state_w_lg_q1765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_data_state_w_lg_q1678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 read_first_nominal_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF read_first_nominal_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_read_first_nominal_state_w_lg_q1773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_first_nominal_state_w_lg_q1684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 read_first_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF read_first_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_read_first_state_w_lg_q1766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_first_state_w_lg_q1676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_first_state_w_lg_w_lg_w_lg_q1894w1895w1896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_first_state_w_lg_w_lg_q1894w1895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_first_state_w_lg_q1894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 read_init_nominal_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF read_init_nominal_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_read_init_nominal_state_w_lg_q1682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 read_init_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF read_init_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_read_init_state_w_lg_q1674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_init_state_w_lg_q1891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 read_last_nominal_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF read_last_nominal_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_read_last_nominal_state_w_lg_q1917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_last_nominal_state_w_lg_q1688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 read_last_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF read_last_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_read_last_state_w_lg_q1680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 reconfig_counter_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reconfig_counter_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_reconfig_counter_state_w_lg_q1700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 reconfig_init_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reconfig_init_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_reconfig_init_state_w_lg_q1698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 reconfig_post_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reconfig_post_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_reconfig_post_state_w_lg_q1849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconfig_post_state_w_lg_q1706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 reconfig_seq_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reconfig_seq_data_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_reconfig_seq_data_state_w_lg_q1704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 reconfig_seq_ena_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reconfig_seq_ena_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_reconfig_seq_ena_state_w_lg_q1903w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_reconfig_seq_ena_state_w_lg_q1904w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_reconfig_seq_ena_state_w_lg_q1702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 reconfig_wait_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reconfig_wait_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_reconfig_wait_state_w_lg_q1853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_reconfig_wait_state_w_lg_q1708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 reset_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '1'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reset_state : SIGNAL IS "POWER_UP_LEVEL=HIGH";

	 SIGNAL  wire_reset_state_w_lg_q1671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rom_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF rom_data_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_rom_data_state_w_lg_q1868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rom_data_state_w_lg_q1889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rom_data_state_w_lg_w_lg_q1897w1933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rom_data_state_w_lg_q1716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rom_data_state_w_lg_w_lg_q1897w1898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rom_data_state_w_lg_w_lg_q1929w1930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rom_data_state_w_lg_q1897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rom_data_state_w_lg_q1929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rom_first_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF rom_first_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_rom_first_state_w_lg_w_lg_w_lg_w_lg_q1943w1944w1945w1947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rom_first_state_w_lg_q1712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rom_first_state_w_lg_w_lg_w_lg_q1943w1944w1945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rom_first_state_w_lg_w_lg_q1943w1944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rom_first_state_w_lg_w_lg_q1885w1886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rom_first_state_w_lg_q1943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rom_first_state_w_lg_q1885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rom_init_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF rom_init_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_rom_init_state_w_lg_q1710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rom_last_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF rom_last_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_rom_last_state_w_lg_q1753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rom_last_state_w_lg_q1720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rom_second_last_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF rom_second_last_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_rom_second_last_state_w_lg_q1754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rom_second_last_state_w_lg_q1718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rom_second_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF rom_second_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_rom_second_state_w_lg_q1714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 shift_reg0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_shift_reg_w_lg_q217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_shift_reg_w_lg_w_lg_q217w218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 shift_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_shift_reg_w_lg_q223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_shift_reg_w_lg_w_lg_q223w224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 shift_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_shift_reg_w_lg_q228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_shift_reg_w_lg_w_lg_q228w229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 shift_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_shift_reg_w_lg_q233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_shift_reg_w_lg_w_lg_q233w234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 shift_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_shift_reg_w_lg_q238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_shift_reg_w_lg_w_lg_q238w239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 shift_reg5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_shift_reg_w_lg_q243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_shift_reg_w_lg_w_lg_q243w244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 shift_reg6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_shift_reg_w_lg_q248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_shift_reg_w_lg_w_lg_q248w249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 shift_reg7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_shift_reg_w_lg_q253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_shift_reg_w_lg_w_lg_q253w254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 shift_reg8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_shift_reg_w_lg_q258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_shift_reg_w_lg_w_lg_q258w259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 shift_reg9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 shift_reg10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 shift_reg11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 shift_reg12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 shift_reg13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 shift_reg14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 shift_reg15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 shift_reg16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 shift_reg17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_shift_reg_w_lg_q262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_shift_reg_w_lg_q264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_shift_reg_w_lg_q267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_shift_reg_w_lg_q270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_shift_reg_w_lg_q273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_shift_reg_w_lg_q276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_shift_reg_w_lg_q279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_shift_reg_w_lg_q282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_shift_reg_ena	:	STD_LOGIC_VECTOR(17 DOWNTO 0);
	 SIGNAL	 tmp_nominal_data_out_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 tmp_seq_ena_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF write_data_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_write_data_state_w_lg_q1738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_data_state_w_lg_q1692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 write_init_nominal_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF write_init_nominal_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_write_init_nominal_state_w_lg_q1694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 write_init_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF write_init_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_write_init_state_w_lg_q1690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_init_state_w_lg_q1900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 write_nominal_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF write_nominal_state : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_write_nominal_state_w_lg_q1737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_nominal_state_w_lg_q1696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_lg_w_result_range214w215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_lg_w_result_range221w222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_lg_w_result_range226w227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_lg_w_result_range231w232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_lg_w_result_range236w237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_lg_w_result_range241w242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_lg_w_result_range246w247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_lg_w_result_range251w252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_lg_w_result_range256w257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_add_sub5_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub5_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub5_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_result_range214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_result_range221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_result_range226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_result_range231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_result_range236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_result_range241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_result_range246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_result_range251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub5_w_result_range256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub6_dataa	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub6_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cmpr7_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr7_dataa	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cmpr7_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cntr1_q	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cntr12_q	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cntr13_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cntr14_q	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cntr15_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_cntr16_q	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cntr2_q	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cntr3_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_decode11_eq	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_addr_counter_out1934w1935w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rom_width_counter_enable1931w1932w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_counter_out1938w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_decoder_out1901w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_c0_wire1828w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_c1_wire1826w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_c2_wire1824w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_c3_wire1822w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_c4_wire1820w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_addr_counter_out1887w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_addr_counter_out1934w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_addr_decoder_out1893w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_reconfig_addr_counter_out1936w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_rom_data_in1946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rom_width_counter_enable1931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rotate_addr_counter_out1937w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_serial_out1948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_counter_param_latch_range294w379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_counter_type_latch_range284w710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dummy_scandataout1925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_pll_scandone1927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_addr_counter_done1867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_nominal_out216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_param1742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reconfig1740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reconfig_done1852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reconfig_post_done1848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reconfig_width_counter_done1845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reset1w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reset_rom_address1752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rom_width_counter_done1888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rotate_width_counter_done1796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_width_counter_done1764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_from_rom1739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_param1741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_counter_param_latch_range296w297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_counter_type_latch_range286w530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w1329w1392w1452w1516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w1329w1392w1452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w1361w1422w1483w1550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w1329w1392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w1361w1422w1483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w1329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w1361w1422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w980w1055w1126w1195w1261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w1361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w980w1055w1126w1195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w1016w1091w1160w1228w1294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w980w1055w1126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w1016w1091w1160w1228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w980w1055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w1016w1091w1160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w1016w1091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w423w570w637w749w817w920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w1016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w423w570w637w749w817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w571w672w784w850w951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_shift_reg_load_enable60w61w62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w423w570w637w749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w571w672w784w850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable60w61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w423w570w637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w571w672w784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dummy_scandataout1926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w301w378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w381w495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w423w570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w571w672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w675w885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  addr_counter_enable :	STD_LOGIC;
	 SIGNAL  addr_counter_out :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  addr_counter_sload :	STD_LOGIC;
	 SIGNAL  addr_counter_sload_value :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  addr_decoder_out :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  c0_wire :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  c1_wire :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  c2_wire :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  c3_wire :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  c4_wire :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  const_scan_chain_size :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  counter_param_latch :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  counter_type_latch :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  cuda_combout_wire :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  dummy_scandataout :	STD_LOGIC;
	 SIGNAL  encode_out :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  input_latch_enable :	STD_LOGIC;
	 SIGNAL  power_up :	STD_LOGIC;
	 SIGNAL  read_addr_counter_done :	STD_LOGIC;
	 SIGNAL  read_addr_counter_enable :	STD_LOGIC;
	 SIGNAL  read_addr_counter_out :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_addr_counter_sload :	STD_LOGIC;
	 SIGNAL  read_addr_counter_sload_value :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_addr_decoder_out :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_nominal_out :	STD_LOGIC;
	 SIGNAL  reconfig_addr_counter_enable :	STD_LOGIC;
	 SIGNAL  reconfig_addr_counter_out :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  reconfig_addr_counter_sload :	STD_LOGIC;
	 SIGNAL  reconfig_addr_counter_sload_value :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  reconfig_done :	STD_LOGIC;
	 SIGNAL  reconfig_post_done :	STD_LOGIC;
	 SIGNAL  reconfig_width_counter_done :	STD_LOGIC;
	 SIGNAL  reconfig_width_counter_enable :	STD_LOGIC;
	 SIGNAL  reconfig_width_counter_sload :	STD_LOGIC;
	 SIGNAL  reconfig_width_counter_sload_value :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  rom_width_counter_done :	STD_LOGIC;
	 SIGNAL  rom_width_counter_enable :	STD_LOGIC;
	 SIGNAL  rom_width_counter_sload :	STD_LOGIC;
	 SIGNAL  rom_width_counter_sload_value :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rotate_addr_counter_enable :	STD_LOGIC;
	 SIGNAL  rotate_addr_counter_out :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rotate_addr_counter_sload :	STD_LOGIC;
	 SIGNAL  rotate_addr_counter_sload_value :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rotate_decoder_wires :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  rotate_width_counter_done :	STD_LOGIC;
	 SIGNAL  rotate_width_counter_enable :	STD_LOGIC;
	 SIGNAL  rotate_width_counter_sload :	STD_LOGIC;
	 SIGNAL  rotate_width_counter_sload_value :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  scan_cache_address :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  scan_cache_in :	STD_LOGIC;
	 SIGNAL  scan_cache_out :	STD_LOGIC;
	 SIGNAL  scan_cache_write_enable :	STD_LOGIC;
	 SIGNAL  sel_param_bypass_LF_unused :	STD_LOGIC;
	 SIGNAL  sel_param_c :	STD_LOGIC;
	 SIGNAL  sel_param_high_i_postscale :	STD_LOGIC;
	 SIGNAL  sel_param_low_r :	STD_LOGIC;
	 SIGNAL  sel_param_nominal_count :	STD_LOGIC;
	 SIGNAL  sel_param_odd_CP_unused :	STD_LOGIC;
	 SIGNAL  sel_type_c0 :	STD_LOGIC;
	 SIGNAL  sel_type_c1 :	STD_LOGIC;
	 SIGNAL  sel_type_c2 :	STD_LOGIC;
	 SIGNAL  sel_type_c3 :	STD_LOGIC;
	 SIGNAL  sel_type_c4 :	STD_LOGIC;
	 SIGNAL  sel_type_cplf :	STD_LOGIC;
	 SIGNAL  sel_type_m :	STD_LOGIC;
	 SIGNAL  sel_type_n :	STD_LOGIC;
	 SIGNAL  sel_type_vco :	STD_LOGIC;
	 SIGNAL  seq_addr_wire :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  seq_sload_value :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  shift_reg_clear :	STD_LOGIC;
	 SIGNAL  shift_reg_load_enable :	STD_LOGIC;
	 SIGNAL  shift_reg_load_nominal_enable :	STD_LOGIC;
	 SIGNAL  shift_reg_serial_in :	STD_LOGIC;
	 SIGNAL  shift_reg_serial_out :	STD_LOGIC;
	 SIGNAL  shift_reg_shift_enable :	STD_LOGIC;
	 SIGNAL  shift_reg_shift_nominal_enable :	STD_LOGIC;
	 SIGNAL  shift_reg_width_select :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  w1019w :	STD_LOGIC;
	 SIGNAL  w1056w :	STD_LOGIC;
	 SIGNAL  w1092w :	STD_LOGIC;
	 SIGNAL  w1127w :	STD_LOGIC;
	 SIGNAL  w1163w :	STD_LOGIC;
	 SIGNAL  w1196w :	STD_LOGIC;
	 SIGNAL  w1229w :	STD_LOGIC;
	 SIGNAL  w1262w :	STD_LOGIC;
	 SIGNAL  w1297w :	STD_LOGIC;
	 SIGNAL  w1330w :	STD_LOGIC;
	 SIGNAL  w1362w :	STD_LOGIC;
	 SIGNAL  w1393w :	STD_LOGIC;
	 SIGNAL  w1424w :	STD_LOGIC;
	 SIGNAL  w1453w :	STD_LOGIC;
	 SIGNAL  w1484w :	STD_LOGIC;
	 SIGNAL  w1517w :	STD_LOGIC;
	 SIGNAL  w1565w :	STD_LOGIC;
	 SIGNAL  w1592w :	STD_LOGIC;
	 SIGNAL  w301w :	STD_LOGIC;
	 SIGNAL  w341w :	STD_LOGIC;
	 SIGNAL  w381w :	STD_LOGIC;
	 SIGNAL  w423w :	STD_LOGIC;
	 SIGNAL  w460w :	STD_LOGIC;
	 SIGNAL  w496w :	STD_LOGIC;
	 SIGNAL  w534w :	STD_LOGIC;
	 SIGNAL  w571w :	STD_LOGIC;
	 SIGNAL  w605w :	STD_LOGIC;
	 SIGNAL  w638w :	STD_LOGIC;
	 SIGNAL  w64w :	STD_LOGIC;
	 SIGNAL  w675w :	STD_LOGIC;
	 SIGNAL  w713w :	STD_LOGIC;
	 SIGNAL  w750w :	STD_LOGIC;
	 SIGNAL  w785w :	STD_LOGIC;
	 SIGNAL  w818w :	STD_LOGIC;
	 SIGNAL  w851w :	STD_LOGIC;
	 SIGNAL  w888w :	STD_LOGIC;
	 SIGNAL  w921w :	STD_LOGIC;
	 SIGNAL  w952w :	STD_LOGIC;
	 SIGNAL  w981w :	STD_LOGIC;
	 SIGNAL  width_counter_done :	STD_LOGIC;
	 SIGNAL  width_counter_enable :	STD_LOGIC;
	 SIGNAL  width_counter_sload :	STD_LOGIC;
	 SIGNAL  width_counter_sload_value :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  width_decoder_out :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  width_decoder_select :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_counter_param_latch_range294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_counter_param_latch_range296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_counter_type_latch_range284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_counter_type_latch_range286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rotate_decoder_wires_range1827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rotate_decoder_wires_range1825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rotate_decoder_wires_range1823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rotate_decoder_wires_range1821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rotate_decoder_wires_range1819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_shift_reg_width_select_range261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_shift_reg_width_select_range263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_shift_reg_width_select_range266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_shift_reg_width_select_range269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_shift_reg_width_select_range272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_shift_reg_width_select_range275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_shift_reg_width_select_range278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_shift_reg_width_select_range281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  altsyncram
	 GENERIC 
	 (
		ADDRESS_ACLR_A	:	STRING := "UNUSED";
		ADDRESS_ACLR_B	:	STRING := "NONE";
		ADDRESS_REG_B	:	STRING := "CLOCK1";
		BYTE_SIZE	:	NATURAL := 8;
		BYTEENA_ACLR_A	:	STRING := "UNUSED";
		BYTEENA_ACLR_B	:	STRING := "NONE";
		BYTEENA_REG_B	:	STRING := "CLOCK1";
		CLOCK_ENABLE_CORE_A	:	STRING := "USE_INPUT_CLKEN";
		CLOCK_ENABLE_CORE_B	:	STRING := "USE_INPUT_CLKEN";
		CLOCK_ENABLE_INPUT_A	:	STRING := "NORMAL";
		CLOCK_ENABLE_INPUT_B	:	STRING := "NORMAL";
		CLOCK_ENABLE_OUTPUT_A	:	STRING := "NORMAL";
		CLOCK_ENABLE_OUTPUT_B	:	STRING := "NORMAL";
		ECC_PIPELINE_STAGE_ENABLED	:	STRING := "FALSE";
		ENABLE_ECC	:	STRING := "FALSE";
		IMPLEMENT_IN_LES	:	STRING := "OFF";
		INDATA_ACLR_A	:	STRING := "UNUSED";
		INDATA_ACLR_B	:	STRING := "NONE";
		INDATA_REG_B	:	STRING := "CLOCK1";
		INIT_FILE	:	STRING := "UNUSED";
		INIT_FILE_LAYOUT	:	STRING := "PORT_A";
		MAXIMUM_DEPTH	:	NATURAL := 0;
		NUMWORDS_A	:	NATURAL := 0;
		NUMWORDS_B	:	NATURAL := 0;
		OPERATION_MODE	:	STRING := "BIDIR_DUAL_PORT";
		OUTDATA_ACLR_A	:	STRING := "NONE";
		OUTDATA_ACLR_B	:	STRING := "NONE";
		OUTDATA_REG_A	:	STRING := "UNREGISTERED";
		OUTDATA_REG_B	:	STRING := "UNREGISTERED";
		POWER_UP_UNINITIALIZED	:	STRING := "FALSE";
		RAM_BLOCK_TYPE	:	STRING := "AUTO";
		RDCONTROL_ACLR_B	:	STRING := "NONE";
		RDCONTROL_REG_B	:	STRING := "CLOCK1";
		READ_DURING_WRITE_MODE_MIXED_PORTS	:	STRING := "DONT_CARE";
		read_during_write_mode_port_a	:	STRING := "NEW_DATA_NO_NBE_READ";
		read_during_write_mode_port_b	:	STRING := "NEW_DATA_NO_NBE_READ";
		WIDTH_A	:	NATURAL;
		WIDTH_B	:	NATURAL := 1;
		WIDTH_BYTEENA_A	:	NATURAL := 1;
		WIDTH_BYTEENA_B	:	NATURAL := 1;
		WIDTH_ECCSTATUS	:	NATURAL := 3;
		WIDTHAD_A	:	NATURAL;
		WIDTHAD_B	:	NATURAL := 1;
		WRCONTROL_ACLR_A	:	STRING := "UNUSED";
		WRCONTROL_ACLR_B	:	STRING := "NONE";
		WRCONTROL_WRADDRESS_REG_B	:	STRING := "CLOCK1";
		INTENDED_DEVICE_FAMILY	:	STRING := "Cyclone 10 LP";
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "altsyncram"
	 );
	 PORT
	 ( 
		aclr0	:	IN STD_LOGIC := '0';
		aclr1	:	IN STD_LOGIC := '0';
		address_a	:	IN STD_LOGIC_VECTOR(WIDTHAD_A-1 DOWNTO 0);
		address_b	:	IN STD_LOGIC_VECTOR(WIDTHAD_B-1 DOWNTO 0) := (OTHERS => '1');
		addressstall_a	:	IN STD_LOGIC := '0';
		addressstall_b	:	IN STD_LOGIC := '0';
		byteena_a	:	IN STD_LOGIC_VECTOR(WIDTH_BYTEENA_A-1 DOWNTO 0) := (OTHERS => '1');
		byteena_b	:	IN STD_LOGIC_VECTOR(WIDTH_BYTEENA_B-1 DOWNTO 0) := (OTHERS => '1');
		clock0	:	IN STD_LOGIC := '1';
		clock1	:	IN STD_LOGIC := '1';
		clocken0	:	IN STD_LOGIC := '1';
		clocken1	:	IN STD_LOGIC := '1';
		clocken2	:	IN STD_LOGIC := '1';
		clocken3	:	IN STD_LOGIC := '1';
		data_a	:	IN STD_LOGIC_VECTOR(WIDTH_A-1 DOWNTO 0) := (OTHERS => '1');
		data_b	:	IN STD_LOGIC_VECTOR(WIDTH_B-1 DOWNTO 0) := (OTHERS => '1');
		eccstatus	:	OUT STD_LOGIC_VECTOR(WIDTH_ECCSTATUS-1 DOWNTO 0);
		q_a	:	OUT STD_LOGIC_VECTOR(WIDTH_A-1 DOWNTO 0);
		q_b	:	OUT STD_LOGIC_VECTOR(WIDTH_B-1 DOWNTO 0);
		rden_a	:	IN STD_LOGIC := '1';
		rden_b	:	IN STD_LOGIC := '1';
		wren_a	:	IN STD_LOGIC := '0';
		wren_b	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  cyclone10lp_lcell_comb
	 GENERIC 
	 (
		DONT_TOUCH	:	STRING := "off";
		LUT_MASK	:	STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000";
		SUM_LUTC_INPUT	:	STRING := "datac";
		lpm_type	:	STRING := "cyclone10lp_lcell_comb"
	 );
	 PORT
	 ( 
		cin	:	IN STD_LOGIC := '0';
		combout	:	OUT STD_LOGIC;
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC := '0';
		datab	:	IN STD_LOGIC := '0';
		datac	:	IN STD_LOGIC := '0';
		datad	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_decode
	 GENERIC 
	 (
		LPM_DECODES	:	NATURAL;
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_decode"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		enable	:	IN STD_LOGIC := '1';
		eq	:	OUT STD_LOGIC_VECTOR(LPM_DECODES-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	loop0 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_read_addr_counter_out1934w1935w(i) <= wire_w_lg_read_addr_counter_out1934w(i) AND wire_rom_data_state_w_lg_w_lg_q1897w1933w(0);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_rom_width_counter_enable1931w1932w(i) <= wire_w_lg_rom_width_counter_enable1931w(0) AND addr_from_rom2(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_addr_counter_out1938w(i) <= addr_counter_out(i) AND addr_counter_enable;
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_addr_decoder_out1901w(i) <= addr_decoder_out(i) AND wire_write_init_state_w_lg_q1900w(0);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_c0_wire1828w(i) <= c0_wire(i) AND wire_w_rotate_decoder_wires_range1827w(0);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_c1_wire1826w(i) <= c1_wire(i) AND wire_w_rotate_decoder_wires_range1825w(0);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_c2_wire1824w(i) <= c2_wire(i) AND wire_w_rotate_decoder_wires_range1823w(0);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_c3_wire1822w(i) <= c3_wire(i) AND wire_w_rotate_decoder_wires_range1821w(0);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_c4_wire1820w(i) <= c4_wire(i) AND wire_w_rotate_decoder_wires_range1819w(0);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_read_addr_counter_out1887w(i) <= read_addr_counter_out(i) AND wire_rom_first_state_w_lg_w_lg_q1885w1886w(0);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_read_addr_counter_out1934w(i) <= read_addr_counter_out(i) AND read_addr_counter_enable;
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_read_addr_decoder_out1893w(i) <= read_addr_decoder_out(i) AND wire_read_init_state_w_lg_q1891w(0);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_reconfig_addr_counter_out1936w(i) <= reconfig_addr_counter_out(i) AND reconfig_addr_counter_enable;
	END GENERATE loop12;
	wire_w_lg_rom_data_in1946w(0) <= rom_data_in AND wire_rom_first_state_w_lg_w_lg_w_lg_q1943w1944w1945w(0);
	wire_w_lg_rom_width_counter_enable1931w(0) <= rom_width_counter_enable AND wire_rom_data_state_w_lg_w_lg_q1929w1930w(0);
	loop13 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_rotate_addr_counter_out1937w(i) <= rotate_addr_counter_out(i) AND rotate_addr_counter_enable;
	END GENERATE loop13;
	wire_w_lg_shift_reg_load_enable187w(0) <= shift_reg_load_enable AND wire_w_data_in_range186w(0);
	wire_w_lg_shift_reg_load_enable179w(0) <= shift_reg_load_enable AND wire_w_data_in_range178w(0);
	wire_w_lg_shift_reg_load_enable171w(0) <= shift_reg_load_enable AND wire_w_data_in_range170w(0);
	wire_w_lg_shift_reg_load_enable163w(0) <= shift_reg_load_enable AND wire_w_data_in_range162w(0);
	wire_w_lg_shift_reg_load_enable155w(0) <= shift_reg_load_enable AND wire_w_data_in_range154w(0);
	wire_w_lg_shift_reg_load_enable147w(0) <= shift_reg_load_enable AND wire_w_data_in_range146w(0);
	wire_w_lg_shift_reg_load_enable139w(0) <= shift_reg_load_enable AND wire_w_data_in_range138w(0);
	wire_w_lg_shift_reg_load_enable131w(0) <= shift_reg_load_enable AND wire_w_data_in_range130w(0);
	wire_w_lg_shift_reg_load_enable123w(0) <= shift_reg_load_enable AND wire_w_data_in_range122w(0);
	wire_w_lg_shift_reg_serial_out1948w(0) <= shift_reg_serial_out AND wire_rom_first_state_w_lg_w_lg_w_lg_w_lg_q1943w1944w1945w1947w(0);
	wire_w_lg_w_counter_param_latch_range294w379w(0) <= wire_w_counter_param_latch_range294w(0) AND wire_w_lg_w_counter_param_latch_range296w297w(0);
	wire_w_lg_w_counter_type_latch_range284w710w(0) <= wire_w_counter_type_latch_range284w(0) AND wire_w_lg_w_counter_type_latch_range286w530w(0);
	wire_w_lg_dummy_scandataout1925w(0) <= NOT dummy_scandataout;
	wire_w_lg_pll_scandone1927w(0) <= NOT pll_scandone;
	wire_w_lg_read_addr_counter_done1867w(0) <= NOT read_addr_counter_done;
	wire_w_lg_read_nominal_out216w(0) <= NOT read_nominal_out;
	wire_w_lg_read_param1742w(0) <= NOT read_param;
	wire_w_lg_reconfig1740w(0) <= NOT reconfig;
	wire_w_lg_reconfig_done1852w(0) <= NOT reconfig_done;
	wire_w_lg_reconfig_post_done1848w(0) <= NOT reconfig_post_done;
	wire_w_lg_reconfig_width_counter_done1845w(0) <= NOT reconfig_width_counter_done;
	wire_w_lg_reset1w(0) <= NOT reset;
	wire_w_lg_reset_rom_address1752w(0) <= NOT reset_rom_address;
	wire_w_lg_rom_width_counter_done1888w(0) <= NOT rom_width_counter_done;
	wire_w_lg_rotate_width_counter_done1796w(0) <= NOT rotate_width_counter_done;
	wire_w_lg_width_counter_done1764w(0) <= NOT width_counter_done;
	wire_w_lg_write_from_rom1739w(0) <= NOT write_from_rom;
	wire_w_lg_write_param1741w(0) <= NOT write_param;
	wire_w_lg_w_counter_param_latch_range296w297w(0) <= NOT wire_w_counter_param_latch_range296w(0);
	wire_w_lg_w_counter_type_latch_range286w530w(0) <= NOT wire_w_counter_type_latch_range286w(0);
	wire_w_lg_w_lg_w_lg_w1329w1392w1452w1516w(0) <= wire_w_lg_w_lg_w1329w1392w1452w(0) OR w1484w;
	wire_w_lg_w_lg_w1329w1392w1452w(0) <= wire_w_lg_w1329w1392w(0) OR w1424w;
	wire_w_lg_w_lg_w_lg_w1361w1422w1483w1550w(0) <= wire_w_lg_w_lg_w1361w1422w1483w(0) OR w1517w;
	wire_w_lg_w1329w1392w(0) <= wire_w1329w(0) OR w1362w;
	wire_w_lg_w_lg_w1361w1422w1483w(0) <= wire_w_lg_w1361w1422w(0) OR w1453w;
	wire_w1329w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w980w1055w1126w1195w1261w(0) OR w1297w;
	wire_w_lg_w1361w1422w(0) <= wire_w1361w(0) OR w1393w;
	wire_w_lg_w_lg_w_lg_w_lg_w980w1055w1126w1195w1261w(0) <= wire_w_lg_w_lg_w_lg_w980w1055w1126w1195w(0) OR w1229w;
	wire_w1361w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w1016w1091w1160w1228w1294w(0) OR w1330w;
	wire_w_lg_w_lg_w_lg_w980w1055w1126w1195w(0) <= wire_w_lg_w_lg_w980w1055w1126w(0) OR w1163w;
	wire_w_lg_w_lg_w_lg_w_lg_w1016w1091w1160w1228w1294w(0) <= wire_w_lg_w_lg_w_lg_w1016w1091w1160w1228w(0) OR w1262w;
	wire_w_lg_w_lg_w980w1055w1126w(0) <= wire_w_lg_w980w1055w(0) OR w1092w;
	wire_w_lg_w_lg_w_lg_w1016w1091w1160w1228w(0) <= wire_w_lg_w_lg_w1016w1091w1160w(0) OR w1196w;
	wire_w_lg_w980w1055w(0) <= wire_w980w(0) OR w1019w;
	wire_w_lg_w_lg_w1016w1091w1160w(0) <= wire_w_lg_w1016w1091w(0) OR w1127w;
	wire_w980w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w423w570w637w749w817w920w(0) OR w952w;
	wire_w_lg_w1016w1091w(0) <= wire_w1016w(0) OR w1056w;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w423w570w637w749w817w920w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w423w570w637w749w817w(0) OR w888w;
	wire_w1016w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w571w672w784w850w951w(0) OR w981w;
	wire_w63w(0) <= wire_w_lg_w_lg_w_lg_shift_reg_load_enable60w61w62w(0) OR shift_reg_clear;
	wire_w_lg_w_lg_w_lg_w_lg_w423w570w637w749w817w(0) <= wire_w_lg_w_lg_w_lg_w423w570w637w749w(0) OR w785w;
	wire_w_lg_w_lg_w_lg_w_lg_w571w672w784w850w951w(0) <= wire_w_lg_w_lg_w_lg_w571w672w784w850w(0) OR w921w;
	wire_w_lg_w_lg_w_lg_shift_reg_load_enable60w61w62w(0) <= wire_w_lg_w_lg_shift_reg_load_enable60w61w(0) OR shift_reg_shift_nominal_enable;
	wire_w_lg_w_lg_w_lg_w423w570w637w749w(0) <= wire_w_lg_w_lg_w423w570w637w(0) OR w713w;
	wire_w_lg_w_lg_w_lg_w571w672w784w850w(0) <= wire_w_lg_w_lg_w571w672w784w(0) OR w818w;
	wire_w_lg_w_lg_shift_reg_load_enable60w61w(0) <= wire_w_lg_shift_reg_load_enable60w(0) OR shift_reg_load_nominal_enable;
	wire_w_lg_w_lg_w423w570w637w(0) <= wire_w_lg_w423w570w(0) OR w605w;
	wire_w_lg_w_lg_w571w672w784w(0) <= wire_w_lg_w571w672w(0) OR w750w;
	wire_w_lg_dummy_scandataout1926w(0) <= dummy_scandataout OR wire_w_lg_dummy_scandataout1925w(0);
	wire_w_lg_shift_reg_load_enable60w(0) <= shift_reg_load_enable OR shift_reg_shift_enable;
	wire_w_lg_w301w378w(0) <= w301w OR w341w;
	wire_w_lg_w381w495w(0) <= w381w OR w460w;
	wire_w_lg_w423w570w(0) <= w423w OR w534w;
	wire_w_lg_w571w672w(0) <= w571w OR w638w;
	wire_w_lg_w675w885w(0) <= w675w OR w851w;
	addr_counter_enable <= (write_data_state OR write_nominal_state);
	addr_counter_out <= wire_cntr1_q;
	addr_counter_sload <= wire_write_init_state_w_lg_q1900w(0);
	addr_counter_sload_value <= wire_w_lg_addr_decoder_out1901w;
	addr_decoder_out <= (((((((((((((((((((((((((((((((((((( "0" & "0" & "0" & "0" & "0" & "0" & "0" & w301w) OR ( "0" & "0" & "0" & "0" & "0" & "0" & w341w & w341w)) OR ( "0" & "0" & "0" & "0" & w381w & "0" & "0" & "0")) OR ( "0" & "0" & "0" & "0" & w423w & "0" & "0" & w423w)) OR ( "0" & "0" & "0" & "0" & w460w & w460w & w460w & "0")) OR ( "0" & "0" & "0" & w496w & "0" & "0" & "0" & w496w)) OR ( "0" & "0" & "0" & w534w & "0" & "0" & w534w & "0")) OR ( "0" & "0" & "0" & w571w & w571w & "0" & w571w & "0")) OR ( "0" & "0" & "0" & w605w & w605w & "0" & w605w & w605w)) OR ( "0" & "0" & w638w & "0" & "0" & "0" & w638w & w638w)) OR ( "0" & "0" & w675w & "0" & "0" & "0" & w675w & w675w)) OR ( "0" & "0" & w713w & "0" & "0" & w713w & "0" & "0")) OR ( "0" & "0" & w750w & "0" & w750w & w750w & "0" & "0")) OR ( "0" & "0" & w785w & "0" & w785w & w785w & "0" & w785w)) OR ( "0" & "0" & w818w & w818w & "0" & w818w & "0" & w818w)) OR ( "0" & "0" & w851w & w851w & "0" & w851w & "0" & w851w)) OR ( "0" & "0" & w888w & w888w & "0" & w888w & w888w & "0")) OR ( "0" & "0" & w921w & w921w & w921w & w921w & w921w & "0")) OR ( "0" & "0" & w952w & w952w & w952w & w952w & w952w & w952w)) OR ( "0" & w981w & "0" & "0" & "0" & w981w & w981w & w981w)) OR ( "0" & w1019w & "0" & "0" & w1019w & "0" & "0" & "0")) OR ( "0" & w1056w & "0" & w1056w & "0" & "0" & "0" & "0")) OR ( "0" & w1092w & "0" & w1092w & "0" & "0" & "0" & w1092w)) OR ( "0" & w1127w & "0" & w1127w & w1127w & "0" & "0" & w1127w)) OR ( "0" & w1163w & "0" & w1163w & w1163w & "0" & w1163w & "0")) OR ( "0" & w1196w & w1196w & "0" & "0" & "0" & w1196w & "0")) OR ( "0" & w1229w & w1229w & "0" & "0" & "0" & w1229w & w1229w)) OR ( "0" & w1262w & w1262w & "0" & w1262w & "0" & w1262w & w1262w)) OR ( "0" & w1297w & w1297w & "0" & w1297w & w1297w & "0" & "0")) OR ( "0" & w1330w & w1330w & w1330w & "0" & w1330w & "0" & "0")) OR ( "0" & w1362w & w1362w & w1362w & "0" & w1362w & "0" & w1362w)) OR ( "0" & w1393w & w1393w & w1393w & w1393w & w1393w & "0" & w1393w)) OR ( "0" & w1424w & w1424w & w1424w & w1424w
 & w1424w & w1424w & "0")) OR ( w1453w & "0" & "0" & "0" & "0" & w1453w & w1453w & "0")) OR ( w1484w & "0" & "0" & "0" & "0" & w1484w & w1484w & w1484w)) OR ( w1517w & "0" & "0" & "0" & w1517w & w1517w & w1517w & w1517w));
	busy <= (wire_idle_state_w_lg_q1672w(0) OR areset_state);
	c0_wire <= "01000111";
	c1_wire <= "01011001";
	c2_wire <= "01101011";
	c3_wire <= "01111101";
	c4_wire <= "10001111";
	const_scan_chain_size <= "10001111";
	counter_param_latch <= counter_param_latch_reg;
	counter_type_latch <= counter_type_latch_reg;
	cuda_combout_wire <= ( wire_le_comb10_combout & wire_le_comb9_combout & wire_le_comb8_combout);
	data_out <= ( wire_shift_reg_w_lg_w_lg_q258w259w & wire_shift_reg_w_lg_w_lg_q253w254w & wire_shift_reg_w_lg_w_lg_q248w249w & wire_shift_reg_w_lg_w_lg_q243w244w & wire_shift_reg_w_lg_w_lg_q238w239w & wire_shift_reg_w_lg_w_lg_q233w234w & wire_shift_reg_w_lg_w_lg_q228w229w & wire_shift_reg_w_lg_w_lg_q223w224w & wire_shift_reg_w_lg_w_lg_q217w218w);
	dummy_scandataout <= pll_scandataout;
	encode_out <= ( C4_ena_state & wire_C2_ena_state_w_lg_q1787w & wire_C1_ena_state_w_lg_q1786w);
	input_latch_enable <= (idle_state AND (write_param OR read_param));
	pll_areset <= (pll_areset_in OR (areset_state AND reconfig_wait_state));
	pll_configupdate <= (configupdate_state AND wire_configupdate3_state_w_lg_q1879w(0));
	pll_scanclk <= clock;
	pll_scanclkena <= ((rotate_width_counter_enable AND wire_w_lg_rotate_width_counter_done1796w(0)) OR reconfig_seq_data_state);
	pll_scandata <= (scan_cache_out AND ((rotate_width_counter_enable OR reconfig_seq_data_state) OR reconfig_post_state));
	power_up <= (((((((((((((((((((((((((wire_reset_state_w_lg_q1671w(0) AND wire_idle_state_w_lg_q1672w(0)) AND wire_read_init_state_w_lg_q1674w(0)) AND wire_read_first_state_w_lg_q1676w(0)) AND wire_read_data_state_w_lg_q1678w(0)) AND wire_read_last_state_w_lg_q1680w(0)) AND wire_read_init_nominal_state_w_lg_q1682w(0)) AND wire_read_first_nominal_state_w_lg_q1684w(0)) AND wire_read_data_nominal_state_w_lg_q1686w(0)) AND wire_read_last_nominal_state_w_lg_q1688w(0)) AND wire_write_init_state_w_lg_q1690w(0)) AND wire_write_data_state_w_lg_q1692w(0)) AND wire_write_init_nominal_state_w_lg_q1694w(0)) AND wire_write_nominal_state_w_lg_q1696w(0)) AND wire_reconfig_init_state_w_lg_q1698w(0)) AND wire_reconfig_counter_state_w_lg_q1700w(0)) AND wire_reconfig_seq_ena_state_w_lg_q1702w(0)) AND wire_reconfig_seq_data_state_w_lg_q1704w(0)) AND wire_reconfig_post_state_w_lg_q1706w(0)) AND wire_reconfig_wait_state_w_lg_q1708w(0)) AND wire_rom_init_state_w_lg_q1710w(0)) AND wire_rom_first_state_w_lg_q1712w(0)) AND wire_rom_second_state_w_lg_q1714w(0)) AND wire_rom_data_state_w_lg_q1716w(0)) AND wire_rom_second_last_state_w_lg_q1718w(0)) AND wire_rom_last_state_w_lg_q1720w(0));
	read_addr_counter_done <= (((((((wire_cntr2_q(0) AND wire_cntr2_q(1)) AND wire_cntr2_q(2)) AND wire_cntr2_q(3)) AND (NOT wire_cntr2_q(4))) AND (NOT wire_cntr2_q(5))) AND (NOT wire_cntr2_q(6))) AND wire_cntr2_q(7));
	read_addr_counter_enable <= (wire_read_first_state_w_lg_w_lg_w_lg_q1894w1895w1896w(0) OR wire_rom_data_state_w_lg_w_lg_q1897w1898w(0));
	read_addr_counter_out <= wire_cntr2_q;
	read_addr_counter_sload <= (wire_read_init_state_w_lg_q1891w(0) OR rom_init_state);
	read_addr_counter_sload_value <= wire_w_lg_read_addr_decoder_out1893w;
	read_addr_decoder_out <= (((((((((((((((((((((((((((((((((((( "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0") OR ( "0" & "0" & "0" & "0" & "0" & "0" & w341w & "0")) OR ( "0" & "0" & "0" & "0" & "0" & w381w & "0" & "0")) OR ( "0" & "0" & "0" & "0" & w423w & "0" & "0" & w423w)) OR ( "0" & "0" & "0" & "0" & w460w & "0" & w460w & "0")) OR ( "0" & "0" & "0" & "0" & w496w & w496w & w496w & w496w)) OR ( "0" & "0" & "0" & w534w & "0" & "0" & w534w & "0")) OR ( "0" & "0" & "0" & w571w & "0" & "0" & w571w & w571w)) OR ( "0" & "0" & "0" & w605w & w605w & "0" & w605w & w605w)) OR ( "0" & "0" & "0" & w638w & w638w & w638w & "0" & "0")) OR ( "0" & "0" & "0" & w675w & "0" & "0" & w675w & "0")) OR ( "0" & "0" & w713w & "0" & "0" & w713w & "0" & "0")) OR ( "0" & "0" & w750w & "0" & "0" & w750w & "0" & w750w)) OR ( "0" & "0" & w785w & "0" & w785w & w785w & "0" & w785w)) OR ( "0" & "0" & w818w & "0" & w818w & w818w & w818w & "0")) OR ( "0" & "0" & w851w & "0" & "0" & w851w & "0" & "0")) OR ( "0" & "0" & w888w & w888w & "0" & w888w & w888w & "0")) OR ( "0" & "0" & w921w & w921w & "0" & w921w & w921w & w921w)) OR ( "0" & "0" & w952w & w952w & w952w & w952w & w952w & w952w)) OR ( "0" & w981w & "0" & "0" & "0" & "0" & "0" & "0")) OR ( "0" & w1019w & "0" & "0" & w1019w & "0" & "0" & "0")) OR ( "0" & w1056w & "0" & "0" & w1056w & "0" & "0" & w1056w)) OR ( "0" & w1092w & "0" & w1092w & "0" & "0" & "0" & w1092w)) OR ( "0" & w1127w & "0" & w1127w & "0" & "0" & w1127w & "0")) OR ( "0" & w1163w & "0" & w1163w & w1163w & "0" & w1163w & "0")) OR ( "0" & w1196w & "0" & w1196w & w1196w & "0" & w1196w & w1196w)) OR ( "0" & w1229w & w1229w & "0" & "0" & "0" & w1229w & w1229w)) OR ( "0" & w1262w & w1262w & "0" & "0" & w1262w & "0" & "0")) OR ( "0" & w1297w & w1297w & "0" & w1297w & w1297w & "0" & "0")) OR ( "0" & w1330w & w1330w & "0" & w1330w & w1330w & "0" & w1330w)) OR ( "0" & w1362w & w1362w & w1362w & "0" & w1362w & "0" & w1362w)) OR ( "0" & w1393w & w1393w & w1393w & "0" & w1393w & w1393w & "0")) OR ( "0" & w1424w & w1424w & w1424w & w1424w & w1424w
 & w1424w & "0")) OR ( "0" & w1453w & w1453w & w1453w & w1453w & w1453w & w1453w & w1453w)) OR ( w1484w & "0" & "0" & "0" & "0" & w1484w & w1484w & w1484w)) OR ( w1517w & "0" & "0" & "0" & w1517w & "0" & "0" & "0"));
	read_nominal_out <= tmp_nominal_data_out_state;
	reconfig_addr_counter_enable <= reconfig_seq_data_state;
	reconfig_addr_counter_out <= wire_cntr12_q;
	reconfig_addr_counter_sload <= reconfig_seq_ena_state;
	reconfig_addr_counter_sload_value <= wire_reconfig_seq_ena_state_w_lg_q1903w;
	reconfig_done <= (wire_w_lg_pll_scandone1927w(0) AND wire_w_lg_dummy_scandataout1926w(0));
	reconfig_post_done <= pll_scandone;
	reconfig_width_counter_done <= ((((((NOT wire_cntr13_q(0)) AND (NOT wire_cntr13_q(1))) AND (NOT wire_cntr13_q(2))) AND (NOT wire_cntr13_q(3))) AND (NOT wire_cntr13_q(4))) AND (NOT wire_cntr13_q(5)));
	reconfig_width_counter_enable <= reconfig_seq_data_state;
	reconfig_width_counter_sload <= reconfig_seq_ena_state;
	reconfig_width_counter_sload_value <= wire_reconfig_seq_ena_state_w_lg_q1904w;
	rom_address_out <= wire_w_lg_read_addr_counter_out1887w;
	rom_width_counter_done <= ((((((((NOT wire_cntr14_q(0)) AND (NOT wire_cntr14_q(1))) AND (NOT wire_cntr14_q(2))) AND (NOT wire_cntr14_q(3))) AND (NOT wire_cntr14_q(4))) AND (NOT wire_cntr14_q(5))) AND (NOT wire_cntr14_q(6))) AND (NOT wire_cntr14_q(7)));
	rom_width_counter_enable <= ((rom_data_state OR rom_last_state) OR rom_second_last_state);
	rom_width_counter_sload <= rom_init_state;
	rom_width_counter_sload_value <= const_scan_chain_size;
	rotate_addr_counter_enable <= ((((C0_data_state OR C1_data_state) OR C2_data_state) OR C3_data_state) OR C4_data_state);
	rotate_addr_counter_out <= wire_cntr16_q;
	rotate_addr_counter_sload <= ((((C0_ena_state OR C1_ena_state) OR C2_ena_state) OR C3_ena_state) OR C4_ena_state);
	rotate_addr_counter_sload_value <= ((((wire_w_lg_c0_wire1828w OR wire_w_lg_c1_wire1826w) OR wire_w_lg_c2_wire1824w) OR wire_w_lg_c3_wire1822w) OR wire_w_lg_c4_wire1820w);
	rotate_decoder_wires <= wire_decode11_eq;
	rotate_width_counter_done <= (((((NOT wire_cntr15_q(0)) AND (NOT wire_cntr15_q(1))) AND (NOT wire_cntr15_q(2))) AND (NOT wire_cntr15_q(3))) AND (NOT wire_cntr15_q(4)));
	rotate_width_counter_enable <= ((((C0_data_state OR C1_data_state) OR C2_data_state) OR C3_data_state) OR C4_data_state);
	rotate_width_counter_sload <= ((((C0_ena_state OR C1_ena_state) OR C2_ena_state) OR C3_ena_state) OR C4_ena_state);
	rotate_width_counter_sload_value <= "10010";
	scan_cache_address <= ((((wire_w_lg_addr_counter_out1938w OR wire_w_lg_rotate_addr_counter_out1937w) OR wire_w_lg_reconfig_addr_counter_out1936w) OR wire_w_lg_w_lg_read_addr_counter_out1934w1935w) OR wire_w_lg_w_lg_rom_width_counter_enable1931w1932w);
	scan_cache_in <= (wire_w_lg_shift_reg_serial_out1948w(0) OR wire_w_lg_rom_data_in1946w(0));
	scan_cache_out <= wire_altsyncram4_q_a(0);
	scan_cache_write_enable <= ((((write_data_state OR write_nominal_state) OR rom_data_state) OR rom_second_last_state) OR rom_last_state);
	sel_param_bypass_LF_unused <= (((NOT counter_param_latch(0)) AND wire_w_lg_w_counter_param_latch_range296w297w(0)) AND counter_param_latch(2));
	sel_param_c <= (((NOT counter_param_latch(0)) AND counter_param_latch(1)) AND (NOT counter_param_latch(2)));
	sel_param_high_i_postscale <= (((NOT counter_param_latch(0)) AND wire_w_lg_w_counter_param_latch_range296w297w(0)) AND (NOT counter_param_latch(2)));
	sel_param_low_r <= (wire_w_lg_w_counter_param_latch_range294w379w(0) AND (NOT counter_param_latch(2)));
	sel_param_nominal_count <= ((counter_param_latch(0) AND counter_param_latch(1)) AND counter_param_latch(2));
	sel_param_odd_CP_unused <= (wire_w_lg_w_counter_param_latch_range294w379w(0) AND counter_param_latch(2));
	sel_type_c0 <= ((((NOT counter_type_latch(0)) AND wire_w_lg_w_counter_type_latch_range286w530w(0)) AND counter_type_latch(2)) AND (NOT counter_type_latch(3)));
	sel_type_c1 <= ((wire_w_lg_w_counter_type_latch_range284w710w(0) AND counter_type_latch(2)) AND (NOT counter_type_latch(3)));
	sel_type_c2 <= ((((NOT counter_type_latch(0)) AND counter_type_latch(1)) AND counter_type_latch(2)) AND (NOT counter_type_latch(3)));
	sel_type_c3 <= (((counter_type_latch(0) AND counter_type_latch(1)) AND counter_type_latch(2)) AND (NOT counter_type_latch(3)));
	sel_type_c4 <= ((((NOT counter_type_latch(0)) AND wire_w_lg_w_counter_type_latch_range286w530w(0)) AND (NOT counter_type_latch(2))) AND counter_type_latch(3));
	sel_type_cplf <= ((((NOT counter_type_latch(0)) AND counter_type_latch(1)) AND (NOT counter_type_latch(2))) AND (NOT counter_type_latch(3)));
	sel_type_m <= ((wire_w_lg_w_counter_type_latch_range284w710w(0) AND (NOT counter_type_latch(2))) AND (NOT counter_type_latch(3)));
	sel_type_n <= ((((NOT counter_type_latch(0)) AND wire_w_lg_w_counter_type_latch_range286w530w(0)) AND (NOT counter_type_latch(2))) AND (NOT counter_type_latch(3)));
	sel_type_vco <= (((counter_type_latch(0) AND counter_type_latch(1)) AND (NOT counter_type_latch(2))) AND (NOT counter_type_latch(3)));
	seq_addr_wire <= "00110101";
	seq_sload_value <= "110110";
	shift_reg_clear <= wire_read_init_state_w_lg_q1891w(0);
	shift_reg_load_enable <= ((idle_state AND write_param) AND (NOT ((((((NOT counter_type(3)) AND (NOT counter_type(2))) AND (NOT counter_type(1))) AND counter_param(2)) AND counter_param(1)) AND counter_param(0))));
	shift_reg_load_nominal_enable <= ((idle_state AND write_param) AND ((((((NOT counter_type(3)) AND (NOT counter_type(2))) AND (NOT counter_type(1))) AND counter_param(2)) AND counter_param(1)) AND counter_param(0)));
	shift_reg_serial_in <= scan_cache_out;
	shift_reg_serial_out <= (((((((wire_shift_reg_w_lg_q262w(0) OR wire_shift_reg_w_lg_q264w(0)) OR wire_shift_reg_w_lg_q267w(0)) OR wire_shift_reg_w_lg_q270w(0)) OR wire_shift_reg_w_lg_q273w(0)) OR wire_shift_reg_w_lg_q276w(0)) OR wire_shift_reg_w_lg_q279w(0)) OR wire_shift_reg_w_lg_q282w(0));
	shift_reg_shift_enable <= ((read_data_state OR read_last_state) OR write_data_state);
	shift_reg_shift_nominal_enable <= ((read_data_nominal_state OR read_last_nominal_state) OR write_nominal_state);
	shift_reg_width_select <= width_decoder_select;
	w1019w <= (sel_type_c1 AND sel_param_bypass_LF_unused);
	w1056w <= (sel_type_c1 AND sel_param_high_i_postscale);
	w1092w <= (sel_type_c1 AND sel_param_odd_CP_unused);
	w1127w <= (sel_type_c1 AND sel_param_low_r);
	w1163w <= (sel_type_c2 AND sel_param_bypass_LF_unused);
	w1196w <= (sel_type_c2 AND sel_param_high_i_postscale);
	w1229w <= (sel_type_c2 AND sel_param_odd_CP_unused);
	w1262w <= (sel_type_c2 AND sel_param_low_r);
	w1297w <= (sel_type_c3 AND sel_param_bypass_LF_unused);
	w1330w <= (sel_type_c3 AND sel_param_high_i_postscale);
	w1362w <= (sel_type_c3 AND sel_param_odd_CP_unused);
	w1393w <= (sel_type_c3 AND sel_param_low_r);
	w1424w <= (sel_type_c4 AND sel_param_bypass_LF_unused);
	w1453w <= (sel_type_c4 AND sel_param_high_i_postscale);
	w1484w <= (sel_type_c4 AND sel_param_odd_CP_unused);
	w1517w <= (sel_type_c4 AND sel_param_low_r);
	w1565w <= '0';
	w1592w <= '0';
	w301w <= (sel_type_cplf AND sel_param_bypass_LF_unused);
	w341w <= (sel_type_cplf AND sel_param_c);
	w381w <= (sel_type_cplf AND sel_param_low_r);
	w423w <= (sel_type_vco AND sel_param_high_i_postscale);
	w460w <= (sel_type_cplf AND sel_param_odd_CP_unused);
	w496w <= (sel_type_cplf AND sel_param_high_i_postscale);
	w534w <= (sel_type_n AND sel_param_bypass_LF_unused);
	w571w <= (sel_type_n AND sel_param_high_i_postscale);
	w605w <= (sel_type_n AND sel_param_odd_CP_unused);
	w638w <= (sel_type_n AND sel_param_low_r);
	w64w <= '0';
	w675w <= (sel_type_n AND sel_param_nominal_count);
	w713w <= (sel_type_m AND sel_param_bypass_LF_unused);
	w750w <= (sel_type_m AND sel_param_high_i_postscale);
	w785w <= (sel_type_m AND sel_param_odd_CP_unused);
	w818w <= (sel_type_m AND sel_param_low_r);
	w851w <= (sel_type_m AND sel_param_nominal_count);
	w888w <= (sel_type_c0 AND sel_param_bypass_LF_unused);
	w921w <= (sel_type_c0 AND sel_param_high_i_postscale);
	w952w <= (sel_type_c0 AND sel_param_odd_CP_unused);
	w981w <= (sel_type_c0 AND sel_param_low_r);
	width_counter_done <= (((((NOT wire_cntr3_q(0)) AND (NOT wire_cntr3_q(1))) AND (NOT wire_cntr3_q(2))) AND (NOT wire_cntr3_q(3))) AND (NOT wire_cntr3_q(4)));
	width_counter_enable <= (((wire_read_first_state_w_lg_q1894w(0) OR write_data_state) OR read_data_nominal_state) OR write_nominal_state);
	width_counter_sload <= (((read_init_state OR write_init_state) OR read_init_nominal_state) OR write_init_nominal_state);
	width_counter_sload_value <= width_decoder_out;
	width_decoder_out <= (((((( "0" & "0" & "0" & "0" & "0") OR ( width_decoder_select(2) & "0" & "0" & "0" & width_decoder_select(2))) OR ( "0" & "0" & "0" & "0" & width_decoder_select(3))) OR ( "0" & "0" & width_decoder_select(5) & width_decoder_select(5) & width_decoder_select(5))) OR ( "0" & "0" & "0" & width_decoder_select(6) & "0")) OR ( "0" & "0" & width_decoder_select(7) & "0" & "0"));
	width_decoder_select <= ( wire_w_lg_w381w495w & w496w & wire_w_lg_w_lg_w_lg_w1361w1422w1483w1550w & w1592w & wire_w_lg_w301w378w & wire_w_lg_w675w885w & w1565w & wire_w_lg_w_lg_w_lg_w1329w1392w1452w1516w);
	write_rom_ena <= (wire_rom_first_state_w_lg_q1885w(0) OR wire_rom_data_state_w_lg_q1889w(0));
	wire_w_counter_param_latch_range294w(0) <= counter_param_latch(0);
	wire_w_counter_param_latch_range296w(0) <= counter_param_latch(1);
	wire_w_counter_type_latch_range284w(0) <= counter_type_latch(0);
	wire_w_counter_type_latch_range286w(0) <= counter_type_latch(1);
	wire_w_data_in_range186w(0) <= data_in(0);
	wire_w_data_in_range178w(0) <= data_in(1);
	wire_w_data_in_range170w(0) <= data_in(2);
	wire_w_data_in_range162w(0) <= data_in(3);
	wire_w_data_in_range154w(0) <= data_in(4);
	wire_w_data_in_range146w(0) <= data_in(5);
	wire_w_data_in_range138w(0) <= data_in(6);
	wire_w_data_in_range130w(0) <= data_in(7);
	wire_w_data_in_range122w(0) <= data_in(8);
	wire_w_rotate_decoder_wires_range1827w(0) <= rotate_decoder_wires(0);
	wire_w_rotate_decoder_wires_range1825w(0) <= rotate_decoder_wires(1);
	wire_w_rotate_decoder_wires_range1823w(0) <= rotate_decoder_wires(2);
	wire_w_rotate_decoder_wires_range1821w(0) <= rotate_decoder_wires(3);
	wire_w_rotate_decoder_wires_range1819w(0) <= rotate_decoder_wires(4);
	wire_w_shift_reg_width_select_range261w(0) <= shift_reg_width_select(0);
	wire_w_shift_reg_width_select_range263w(0) <= shift_reg_width_select(1);
	wire_w_shift_reg_width_select_range266w(0) <= shift_reg_width_select(2);
	wire_w_shift_reg_width_select_range269w(0) <= shift_reg_width_select(3);
	wire_w_shift_reg_width_select_range272w(0) <= shift_reg_width_select(4);
	wire_w_shift_reg_width_select_range275w(0) <= shift_reg_width_select(5);
	wire_w_shift_reg_width_select_range278w(0) <= shift_reg_width_select(6);
	wire_w_shift_reg_width_select_range281w(0) <= shift_reg_width_select(7);
	wire_altsyncram4_data_a(0) <= ( scan_cache_in);
	altsyncram4 :  altsyncram
	  GENERIC MAP (
		INIT_FILE => "./Atari800XL/mist/ntsc.mif",
		NUMWORDS_A => 144,
		OPERATION_MODE => "SINGLE_PORT",
		WIDTH_A => 1,
		WIDTH_BYTEENA_A => 1,
		WIDTHAD_A => 8,
		INTENDED_DEVICE_FAMILY => "Cyclone 10 LP"
	  )
	  PORT MAP ( 
		address_a => scan_cache_address,
		clock0 => clock,
		data_a => wire_altsyncram4_data_a,
		q_a => wire_altsyncram4_q_a,
		wren_a => scan_cache_write_enable
	  );
	le_comb10 :  cyclone10lp_lcell_comb
	  GENERIC MAP (
		DONT_TOUCH => "on",
		LUT_MASK => "1111000011110000",
		SUM_LUTC_INPUT => "datac"
	  )
	  PORT MAP ( 
		combout => wire_le_comb10_combout,
		dataa => encode_out(0),
		datab => encode_out(1),
		datac => encode_out(2)
	  );
	le_comb8 :  cyclone10lp_lcell_comb
	  GENERIC MAP (
		DONT_TOUCH => "on",
		LUT_MASK => "1010101010101010",
		SUM_LUTC_INPUT => "datac"
	  )
	  PORT MAP ( 
		combout => wire_le_comb8_combout,
		dataa => encode_out(0),
		datab => encode_out(1),
		datac => encode_out(2)
	  );
	le_comb9 :  cyclone10lp_lcell_comb
	  GENERIC MAP (
		DONT_TOUCH => "on",
		LUT_MASK => "1100110011001100",
		SUM_LUTC_INPUT => "datac"
	  )
	  PORT MAP ( 
		combout => wire_le_comb9_combout,
		dataa => encode_out(0),
		datab => encode_out(1),
		datac => encode_out(2)
	  );
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN addr_from_rom <= read_addr_counter_out;
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN addr_from_rom2 <= addr_from_rom;
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN areset_init_state_1 <= pll_scandone;
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN areset_state <= (areset_init_state_1 AND wire_w_lg_reset1w(0));
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN C0_data_state <= (C0_ena_state OR (C0_data_state AND wire_w_lg_rotate_width_counter_done1796w(0)));
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN C0_ena_state <= (C1_data_state AND rotate_width_counter_done);
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN C1_data_state <= (C1_ena_state OR (C1_data_state AND wire_w_lg_rotate_width_counter_done1796w(0)));
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN C1_ena_state <= (C2_data_state AND rotate_width_counter_done);
		END IF;
	END PROCESS;
	wire_C1_ena_state_w_lg_q1786w(0) <= C1_ena_state OR C3_ena_state;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN C2_data_state <= (C2_ena_state OR (C2_data_state AND wire_w_lg_rotate_width_counter_done1796w(0)));
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN C2_ena_state <= (C3_data_state AND rotate_width_counter_done);
		END IF;
	END PROCESS;
	wire_C2_ena_state_w_lg_q1787w(0) <= C2_ena_state OR C3_ena_state;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN C3_data_state <= (C3_ena_state OR (C3_data_state AND wire_w_lg_rotate_width_counter_done1796w(0)));
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN C3_ena_state <= (C4_data_state AND rotate_width_counter_done);
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN C4_data_state <= (C4_ena_state OR (C4_data_state AND wire_w_lg_rotate_width_counter_done1796w(0)));
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN C4_ena_state <= reconfig_init_state;
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN configupdate2_state <= configupdate_state;
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '0' AND clock'event) THEN configupdate3_state <= configupdate2_state;
		END IF;
	END PROCESS;
	wire_configupdate3_state_w_lg_q1879w(0) <= NOT configupdate3_state;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN configupdate_state <= reconfig_post_state;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN counter_param_latch_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (input_latch_enable = '1') THEN counter_param_latch_reg <= counter_param;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN counter_type_latch_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (input_latch_enable = '1') THEN counter_type_latch_reg <= counter_type;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN idle_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN idle_state <= (((((wire_idle_state_w_lg_w_lg_w_lg_w1747w1748w1749w1750w(0) OR (reconfig_wait_state AND reconfig_done)) OR ((rom_data_state AND rom_width_counter_done) AND wire_w_lg_reset_rom_address1752w(0))) OR wire_rom_second_last_state_w_lg_q1754w(0)) OR wire_rom_last_state_w_lg_q1753w(0)) OR reset_state);
		END IF;
	END PROCESS;
	wire_idle_state_w_lg_w_lg_w_lg_w_lg_q1743w1744w1745w1746w(0) <= wire_idle_state_w_lg_w_lg_w_lg_q1743w1744w1745w(0) AND wire_w_lg_write_from_rom1739w(0);
	wire_idle_state_w_lg_w_lg_w_lg_q1743w1744w1745w(0) <= wire_idle_state_w_lg_w_lg_q1743w1744w(0) AND wire_w_lg_reconfig1740w(0);
	wire_idle_state_w_lg_w_lg_q1743w1744w(0) <= wire_idle_state_w_lg_q1743w(0) AND wire_w_lg_write_param1741w(0);
	wire_idle_state_w_lg_q1743w(0) <= idle_state AND wire_w_lg_read_param1742w(0);
	wire_idle_state_w_lg_q1672w(0) <= NOT idle_state;
	wire_idle_state_w1747w(0) <= wire_idle_state_w_lg_w_lg_w_lg_w_lg_q1743w1744w1745w1746w(0) OR read_last_state;
	wire_idle_state_w_lg_w1747w1748w(0) <= wire_idle_state_w1747w(0) OR wire_write_data_state_w_lg_q1738w(0);
	wire_idle_state_w_lg_w_lg_w1747w1748w1749w(0) <= wire_idle_state_w_lg_w1747w1748w(0) OR wire_write_nominal_state_w_lg_q1737w(0);
	wire_idle_state_w_lg_w_lg_w_lg_w1747w1748w1749w1750w(0) <= wire_idle_state_w_lg_w_lg_w1747w1748w1749w(0) OR read_last_nominal_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data0 <= wire_add_sub6_result(0);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data1 <= wire_add_sub6_result(1);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data2 <= wire_add_sub6_result(2);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data3 <= wire_add_sub6_result(3);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data4 <= wire_add_sub6_result(4);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data5 <= wire_add_sub6_result(5);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data6 <= wire_add_sub6_result(6);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data7 <= wire_add_sub6_result(7);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data8 <= wire_w_data_in_range186w(0);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data9 <= wire_w_data_in_range178w(0);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data10 <= wire_w_data_in_range170w(0);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data11 <= wire_w_data_in_range162w(0);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data12 <= wire_w_data_in_range154w(0);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data13 <= wire_w_data_in_range146w(0);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data14 <= wire_w_data_in_range138w(0);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data15 <= wire_w_data_in_range130w(0);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data16 <= wire_w_data_in_range122w(0);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN nominal_data17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN nominal_data17 <= wire_cmpr7_aeb;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_data_nominal_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_data_nominal_state <= (wire_read_first_nominal_state_w_lg_q1773w(0) OR wire_read_data_nominal_state_w_lg_q1772w(0));
		END IF;
	END PROCESS;
	wire_read_data_nominal_state_w_lg_q1772w(0) <= read_data_nominal_state AND wire_w_lg_width_counter_done1764w(0);
	wire_read_data_nominal_state_w_lg_q1686w(0) <= NOT read_data_nominal_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_data_state <= (wire_read_first_state_w_lg_q1766w(0) OR wire_read_data_state_w_lg_q1765w(0));
		END IF;
	END PROCESS;
	wire_read_data_state_w_lg_q1765w(0) <= read_data_state AND wire_w_lg_width_counter_done1764w(0);
	wire_read_data_state_w_lg_q1678w(0) <= NOT read_data_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_first_nominal_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_first_nominal_state <= read_init_nominal_state;
		END IF;
	END PROCESS;
	wire_read_first_nominal_state_w_lg_q1773w(0) <= read_first_nominal_state AND wire_w_lg_width_counter_done1764w(0);
	wire_read_first_nominal_state_w_lg_q1684w(0) <= NOT read_first_nominal_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_first_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_first_state <= read_init_state;
		END IF;
	END PROCESS;
	wire_read_first_state_w_lg_q1766w(0) <= read_first_state AND wire_w_lg_width_counter_done1764w(0);
	wire_read_first_state_w_lg_q1676w(0) <= NOT read_first_state;
	wire_read_first_state_w_lg_w_lg_w_lg_q1894w1895w1896w(0) <= wire_read_first_state_w_lg_w_lg_q1894w1895w(0) OR read_data_nominal_state;
	wire_read_first_state_w_lg_w_lg_q1894w1895w(0) <= wire_read_first_state_w_lg_q1894w(0) OR read_first_nominal_state;
	wire_read_first_state_w_lg_q1894w(0) <= read_first_state OR read_data_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_init_nominal_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_init_nominal_state <= ((idle_state AND read_param) AND ((((((NOT counter_type(3)) AND (NOT counter_type(2))) AND (NOT counter_type(1))) AND counter_param(2)) AND counter_param(1)) AND counter_param(0)));
		END IF;
	END PROCESS;
	wire_read_init_nominal_state_w_lg_q1682w(0) <= NOT read_init_nominal_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_init_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_init_state <= ((idle_state AND read_param) AND (NOT ((((((NOT counter_type(3)) AND (NOT counter_type(2))) AND (NOT counter_type(1))) AND counter_param(2)) AND counter_param(1)) AND counter_param(0))));
		END IF;
	END PROCESS;
	wire_read_init_state_w_lg_q1674w(0) <= NOT read_init_state;
	wire_read_init_state_w_lg_q1891w(0) <= read_init_state OR read_init_nominal_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_last_nominal_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_last_nominal_state <= ((read_first_nominal_state AND width_counter_done) OR (read_data_nominal_state AND width_counter_done));
		END IF;
	END PROCESS;
	wire_read_last_nominal_state_w_lg_q1917w(0) <= read_last_nominal_state AND wire_idle_state_w_lg_q1672w(0);
	wire_read_last_nominal_state_w_lg_q1688w(0) <= NOT read_last_nominal_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_last_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_last_state <= ((read_first_state AND width_counter_done) OR (read_data_state AND width_counter_done));
		END IF;
	END PROCESS;
	wire_read_last_state_w_lg_q1680w(0) <= NOT read_last_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN reconfig_counter_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN reconfig_counter_state <= ((((((((((reconfig_init_state OR C0_data_state) OR C1_data_state) OR C2_data_state) OR C3_data_state) OR C4_data_state) OR C0_ena_state) OR C1_ena_state) OR C2_ena_state) OR C3_ena_state) OR C4_ena_state);
		END IF;
	END PROCESS;
	wire_reconfig_counter_state_w_lg_q1700w(0) <= NOT reconfig_counter_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN reconfig_init_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN reconfig_init_state <= (idle_state AND reconfig);
		END IF;
	END PROCESS;
	wire_reconfig_init_state_w_lg_q1698w(0) <= NOT reconfig_init_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN reconfig_post_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN reconfig_post_state <= ((reconfig_seq_data_state AND reconfig_width_counter_done) OR wire_reconfig_post_state_w_lg_q1849w(0));
		END IF;
	END PROCESS;
	wire_reconfig_post_state_w_lg_q1849w(0) <= reconfig_post_state AND wire_w_lg_reconfig_post_done1848w(0);
	wire_reconfig_post_state_w_lg_q1706w(0) <= NOT reconfig_post_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN reconfig_seq_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN reconfig_seq_data_state <= (reconfig_seq_ena_state OR (reconfig_seq_data_state AND wire_w_lg_reconfig_width_counter_done1845w(0)));
		END IF;
	END PROCESS;
	wire_reconfig_seq_data_state_w_lg_q1704w(0) <= NOT reconfig_seq_data_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN reconfig_seq_ena_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN reconfig_seq_ena_state <= tmp_seq_ena_state;
		END IF;
	END PROCESS;
	loop14 : FOR i IN 0 TO 7 GENERATE 
		wire_reconfig_seq_ena_state_w_lg_q1903w(i) <= reconfig_seq_ena_state AND seq_addr_wire(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 5 GENERATE 
		wire_reconfig_seq_ena_state_w_lg_q1904w(i) <= reconfig_seq_ena_state AND seq_sload_value(i);
	END GENERATE loop15;
	wire_reconfig_seq_ena_state_w_lg_q1702w(0) <= NOT reconfig_seq_ena_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN reconfig_wait_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN reconfig_wait_state <= ((reconfig_post_state AND reconfig_post_done) OR wire_reconfig_wait_state_w_lg_q1853w(0));
		END IF;
	END PROCESS;
	wire_reconfig_wait_state_w_lg_q1853w(0) <= reconfig_wait_state AND wire_w_lg_reconfig_done1852w(0);
	wire_reconfig_wait_state_w_lg_q1708w(0) <= NOT reconfig_wait_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN reset_state <= '1';
		ELSIF (clock = '1' AND clock'event) THEN reset_state <= power_up;
		END IF;
	END PROCESS;
	wire_reset_state_w_lg_q1671w(0) <= NOT reset_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN rom_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN rom_data_state <= (rom_second_state OR (wire_rom_data_state_w_lg_q1868w(0) AND wire_w_lg_reset_rom_address1752w(0)));
		END IF;
	END PROCESS;
	wire_rom_data_state_w_lg_q1868w(0) <= rom_data_state AND wire_w_lg_read_addr_counter_done1867w(0);
	wire_rom_data_state_w_lg_q1889w(0) <= rom_data_state AND wire_w_lg_rom_width_counter_done1888w(0);
	wire_rom_data_state_w_lg_w_lg_q1897w1933w(0) <= NOT wire_rom_data_state_w_lg_q1897w(0);
	wire_rom_data_state_w_lg_q1716w(0) <= NOT rom_data_state;
	wire_rom_data_state_w_lg_w_lg_q1897w1898w(0) <= wire_rom_data_state_w_lg_q1897w(0) OR rom_second_state;
	wire_rom_data_state_w_lg_w_lg_q1929w1930w(0) <= wire_rom_data_state_w_lg_q1929w(0) OR rom_last_state;
	wire_rom_data_state_w_lg_q1897w(0) <= rom_data_state OR rom_first_state;
	wire_rom_data_state_w_lg_q1929w(0) <= rom_data_state OR rom_second_last_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN rom_first_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN rom_first_state <= rom_init_state;
		END IF;
	END PROCESS;
	wire_rom_first_state_w_lg_w_lg_w_lg_w_lg_q1943w1944w1945w1947w(0) <= NOT wire_rom_first_state_w_lg_w_lg_w_lg_q1943w1944w1945w(0);
	wire_rom_first_state_w_lg_q1712w(0) <= NOT rom_first_state;
	wire_rom_first_state_w_lg_w_lg_w_lg_q1943w1944w1945w(0) <= wire_rom_first_state_w_lg_w_lg_q1943w1944w(0) OR rom_last_state;
	wire_rom_first_state_w_lg_w_lg_q1943w1944w(0) <= wire_rom_first_state_w_lg_q1943w(0) OR rom_second_last_state;
	wire_rom_first_state_w_lg_w_lg_q1885w1886w(0) <= wire_rom_first_state_w_lg_q1885w(0) OR rom_data_state;
	wire_rom_first_state_w_lg_q1943w(0) <= rom_first_state OR rom_data_state;
	wire_rom_first_state_w_lg_q1885w(0) <= rom_first_state OR rom_second_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN rom_init_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN rom_init_state <= (((((idle_state AND write_from_rom) OR (rom_first_state AND reset_rom_address)) OR (rom_second_state AND reset_rom_address)) OR (rom_data_state AND reset_rom_address)) OR (rom_second_last_state AND reset_rom_address));
		END IF;
	END PROCESS;
	wire_rom_init_state_w_lg_q1710w(0) <= NOT rom_init_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN rom_last_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN rom_last_state <= wire_rom_second_last_state_w_lg_q1754w(0);
		END IF;
	END PROCESS;
	wire_rom_last_state_w_lg_q1753w(0) <= rom_last_state AND wire_w_lg_reset_rom_address1752w(0);
	wire_rom_last_state_w_lg_q1720w(0) <= NOT rom_last_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN rom_second_last_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN rom_second_last_state <= ((rom_data_state AND read_addr_counter_done) AND wire_w_lg_reset_rom_address1752w(0));
		END IF;
	END PROCESS;
	wire_rom_second_last_state_w_lg_q1754w(0) <= rom_second_last_state AND wire_w_lg_reset_rom_address1752w(0);
	wire_rom_second_last_state_w_lg_q1718w(0) <= NOT rom_second_last_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN rom_second_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN rom_second_state <= (rom_first_state AND wire_w_lg_reset_rom_address1752w(0));
		END IF;
	END PROCESS;
	wire_rom_second_state_w_lg_q1714w(0) <= NOT rom_second_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(0) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg0 <= '0';
				ELSE shift_reg0 <= ((((shift_reg_load_nominal_enable AND nominal_data17) OR (shift_reg_load_enable AND w64w)) OR (shift_reg_shift_enable AND shift_reg_serial_in)) OR (shift_reg_shift_nominal_enable AND shift_reg_serial_in));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_shift_reg_w_lg_q217w(0) <= shift_reg0 AND wire_w_lg_read_nominal_out216w(0);
	wire_shift_reg_w_lg_w_lg_q217w218w(0) <= wire_shift_reg_w_lg_q217w(0) OR wire_add_sub5_w_lg_w_result_range214w215w(0);
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(1) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg1 <= '0';
				ELSE shift_reg1 <= ((((shift_reg_load_nominal_enable AND nominal_data16) OR (shift_reg_load_enable AND w64w)) OR (shift_reg_shift_enable AND shift_reg0)) OR (shift_reg_shift_nominal_enable AND shift_reg0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_shift_reg_w_lg_q223w(0) <= shift_reg1 AND wire_w_lg_read_nominal_out216w(0);
	wire_shift_reg_w_lg_w_lg_q223w224w(0) <= wire_shift_reg_w_lg_q223w(0) OR wire_add_sub5_w_lg_w_result_range221w222w(0);
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(2) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg2 <= '0';
				ELSE shift_reg2 <= ((((shift_reg_load_nominal_enable AND nominal_data15) OR (shift_reg_load_enable AND w64w)) OR (shift_reg_shift_enable AND shift_reg1)) OR (shift_reg_shift_nominal_enable AND shift_reg1));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_shift_reg_w_lg_q228w(0) <= shift_reg2 AND wire_w_lg_read_nominal_out216w(0);
	wire_shift_reg_w_lg_w_lg_q228w229w(0) <= wire_shift_reg_w_lg_q228w(0) OR wire_add_sub5_w_lg_w_result_range226w227w(0);
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(3) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg3 <= '0';
				ELSE shift_reg3 <= ((((shift_reg_load_nominal_enable AND nominal_data14) OR (shift_reg_load_enable AND w64w)) OR (shift_reg_shift_enable AND shift_reg2)) OR (shift_reg_shift_nominal_enable AND shift_reg2));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_shift_reg_w_lg_q233w(0) <= shift_reg3 AND wire_w_lg_read_nominal_out216w(0);
	wire_shift_reg_w_lg_w_lg_q233w234w(0) <= wire_shift_reg_w_lg_q233w(0) OR wire_add_sub5_w_lg_w_result_range231w232w(0);
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(4) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg4 <= '0';
				ELSE shift_reg4 <= ((((shift_reg_load_nominal_enable AND nominal_data13) OR (shift_reg_load_enable AND w64w)) OR (shift_reg_shift_enable AND shift_reg3)) OR (shift_reg_shift_nominal_enable AND shift_reg3));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_shift_reg_w_lg_q238w(0) <= shift_reg4 AND wire_w_lg_read_nominal_out216w(0);
	wire_shift_reg_w_lg_w_lg_q238w239w(0) <= wire_shift_reg_w_lg_q238w(0) OR wire_add_sub5_w_lg_w_result_range236w237w(0);
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(5) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg5 <= '0';
				ELSE shift_reg5 <= ((((shift_reg_load_nominal_enable AND nominal_data12) OR (shift_reg_load_enable AND w64w)) OR (shift_reg_shift_enable AND shift_reg4)) OR (shift_reg_shift_nominal_enable AND shift_reg4));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_shift_reg_w_lg_q243w(0) <= shift_reg5 AND wire_w_lg_read_nominal_out216w(0);
	wire_shift_reg_w_lg_w_lg_q243w244w(0) <= wire_shift_reg_w_lg_q243w(0) OR wire_add_sub5_w_lg_w_result_range241w242w(0);
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(6) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg6 <= '0';
				ELSE shift_reg6 <= ((((shift_reg_load_nominal_enable AND nominal_data11) OR (shift_reg_load_enable AND w64w)) OR (shift_reg_shift_enable AND shift_reg5)) OR (shift_reg_shift_nominal_enable AND shift_reg5));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_shift_reg_w_lg_q248w(0) <= shift_reg6 AND wire_w_lg_read_nominal_out216w(0);
	wire_shift_reg_w_lg_w_lg_q248w249w(0) <= wire_shift_reg_w_lg_q248w(0) OR wire_add_sub5_w_lg_w_result_range246w247w(0);
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(7) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg7 <= '0';
				ELSE shift_reg7 <= ((((shift_reg_load_nominal_enable AND nominal_data10) OR (shift_reg_load_enable AND w64w)) OR (shift_reg_shift_enable AND shift_reg6)) OR (shift_reg_shift_nominal_enable AND shift_reg6));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_shift_reg_w_lg_q253w(0) <= shift_reg7 AND wire_w_lg_read_nominal_out216w(0);
	wire_shift_reg_w_lg_w_lg_q253w254w(0) <= wire_shift_reg_w_lg_q253w(0) OR wire_add_sub5_w_lg_w_result_range251w252w(0);
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(8) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg8 <= '0';
				ELSE shift_reg8 <= ((((shift_reg_load_nominal_enable AND nominal_data9) OR (shift_reg_load_enable AND w64w)) OR (shift_reg_shift_enable AND shift_reg7)) OR (shift_reg_shift_nominal_enable AND shift_reg7));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_shift_reg_w_lg_q258w(0) <= shift_reg8 AND wire_w_lg_read_nominal_out216w(0);
	wire_shift_reg_w_lg_w_lg_q258w259w(0) <= wire_shift_reg_w_lg_q258w(0) OR wire_add_sub5_w_lg_w_result_range256w257w(0);
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(9) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg9 <= '0';
				ELSE shift_reg9 <= ((((shift_reg_load_nominal_enable AND nominal_data8) OR wire_w_lg_shift_reg_load_enable123w(0)) OR (shift_reg_shift_enable AND shift_reg8)) OR (shift_reg_shift_nominal_enable AND shift_reg8));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(10) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg10 <= '0';
				ELSE shift_reg10 <= ((((shift_reg_load_nominal_enable AND nominal_data7) OR wire_w_lg_shift_reg_load_enable131w(0)) OR (shift_reg_shift_enable AND shift_reg9)) OR (shift_reg_shift_nominal_enable AND shift_reg9));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(11) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg11 <= '0';
				ELSE shift_reg11 <= ((((shift_reg_load_nominal_enable AND nominal_data6) OR wire_w_lg_shift_reg_load_enable139w(0)) OR (shift_reg_shift_enable AND shift_reg10)) OR (shift_reg_shift_nominal_enable AND shift_reg10));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(12) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg12 <= '0';
				ELSE shift_reg12 <= ((((shift_reg_load_nominal_enable AND nominal_data5) OR wire_w_lg_shift_reg_load_enable147w(0)) OR (shift_reg_shift_enable AND shift_reg11)) OR (shift_reg_shift_nominal_enable AND shift_reg11));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(13) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg13 <= '0';
				ELSE shift_reg13 <= ((((shift_reg_load_nominal_enable AND nominal_data4) OR wire_w_lg_shift_reg_load_enable155w(0)) OR (shift_reg_shift_enable AND shift_reg12)) OR (shift_reg_shift_nominal_enable AND shift_reg12));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(14) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg14 <= '0';
				ELSE shift_reg14 <= ((((shift_reg_load_nominal_enable AND nominal_data3) OR wire_w_lg_shift_reg_load_enable163w(0)) OR (shift_reg_shift_enable AND shift_reg13)) OR (shift_reg_shift_nominal_enable AND shift_reg13));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(15) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg15 <= '0';
				ELSE shift_reg15 <= ((((shift_reg_load_nominal_enable AND nominal_data2) OR wire_w_lg_shift_reg_load_enable171w(0)) OR (shift_reg_shift_enable AND shift_reg14)) OR (shift_reg_shift_nominal_enable AND shift_reg14));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(16) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg16 <= '0';
				ELSE shift_reg16 <= ((((shift_reg_load_nominal_enable AND nominal_data1) OR wire_w_lg_shift_reg_load_enable179w(0)) OR (shift_reg_shift_enable AND shift_reg15)) OR (shift_reg_shift_nominal_enable AND shift_reg15));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN shift_reg17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_shift_reg_ena(17) = '1') THEN 
				IF (shift_reg_clear = '1') THEN shift_reg17 <= '0';
				ELSE shift_reg17 <= ((((shift_reg_load_nominal_enable AND nominal_data0) OR wire_w_lg_shift_reg_load_enable187w(0)) OR (shift_reg_shift_enable AND shift_reg16)) OR (shift_reg_shift_nominal_enable AND shift_reg16));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_shift_reg_w_lg_q262w(0) <= shift_reg17 AND wire_w_shift_reg_width_select_range261w(0);
	wire_shift_reg_w_lg_q264w(0) <= shift_reg17 AND wire_w_shift_reg_width_select_range263w(0);
	wire_shift_reg_w_lg_q267w(0) <= shift_reg17 AND wire_w_shift_reg_width_select_range266w(0);
	wire_shift_reg_w_lg_q270w(0) <= shift_reg17 AND wire_w_shift_reg_width_select_range269w(0);
	wire_shift_reg_w_lg_q273w(0) <= shift_reg17 AND wire_w_shift_reg_width_select_range272w(0);
	wire_shift_reg_w_lg_q276w(0) <= shift_reg17 AND wire_w_shift_reg_width_select_range275w(0);
	wire_shift_reg_w_lg_q279w(0) <= shift_reg17 AND wire_w_shift_reg_width_select_range278w(0);
	wire_shift_reg_w_lg_q282w(0) <= shift_reg17 AND wire_w_shift_reg_width_select_range281w(0);
	loop16 : FOR i IN 0 TO 17 GENERATE
		wire_shift_reg_ena(i) <= wire_w63w(0);
	END GENERATE loop16;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN tmp_nominal_data_out_state <= (wire_read_last_nominal_state_w_lg_q1917w(0) OR (tmp_nominal_data_out_state AND idle_state));
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN tmp_seq_ena_state <= (reconfig_counter_state AND (C0_data_state AND rotate_width_counter_done));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_data_state <= (write_init_state OR (write_data_state AND wire_w_lg_width_counter_done1764w(0)));
		END IF;
	END PROCESS;
	wire_write_data_state_w_lg_q1738w(0) <= write_data_state AND width_counter_done;
	wire_write_data_state_w_lg_q1692w(0) <= NOT write_data_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_init_nominal_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_init_nominal_state <= ((idle_state AND write_param) AND ((((((NOT counter_type(3)) AND (NOT counter_type(2))) AND (NOT counter_type(1))) AND counter_param(2)) AND counter_param(1)) AND counter_param(0)));
		END IF;
	END PROCESS;
	wire_write_init_nominal_state_w_lg_q1694w(0) <= NOT write_init_nominal_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_init_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_init_state <= ((idle_state AND write_param) AND (NOT ((((((NOT counter_type(3)) AND (NOT counter_type(2))) AND (NOT counter_type(1))) AND counter_param(2)) AND counter_param(1)) AND counter_param(0))));
		END IF;
	END PROCESS;
	wire_write_init_state_w_lg_q1690w(0) <= NOT write_init_state;
	wire_write_init_state_w_lg_q1900w(0) <= write_init_state OR write_init_nominal_state;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_nominal_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_nominal_state <= (write_init_nominal_state OR (write_nominal_state AND wire_w_lg_width_counter_done1764w(0)));
		END IF;
	END PROCESS;
	wire_write_nominal_state_w_lg_q1737w(0) <= write_nominal_state AND width_counter_done;
	wire_write_nominal_state_w_lg_q1696w(0) <= NOT write_nominal_state;
	wire_add_sub5_w_lg_w_result_range214w215w(0) <= wire_add_sub5_w_result_range214w(0) AND read_nominal_out;
	wire_add_sub5_w_lg_w_result_range221w222w(0) <= wire_add_sub5_w_result_range221w(0) AND read_nominal_out;
	wire_add_sub5_w_lg_w_result_range226w227w(0) <= wire_add_sub5_w_result_range226w(0) AND read_nominal_out;
	wire_add_sub5_w_lg_w_result_range231w232w(0) <= wire_add_sub5_w_result_range231w(0) AND read_nominal_out;
	wire_add_sub5_w_lg_w_result_range236w237w(0) <= wire_add_sub5_w_result_range236w(0) AND read_nominal_out;
	wire_add_sub5_w_lg_w_result_range241w242w(0) <= wire_add_sub5_w_result_range241w(0) AND read_nominal_out;
	wire_add_sub5_w_lg_w_result_range246w247w(0) <= wire_add_sub5_w_result_range246w(0) AND read_nominal_out;
	wire_add_sub5_w_lg_w_result_range251w252w(0) <= wire_add_sub5_w_result_range251w(0) AND read_nominal_out;
	wire_add_sub5_w_lg_w_result_range256w257w(0) <= wire_add_sub5_w_result_range256w(0) AND read_nominal_out;
	wire_add_sub5_dataa <= ( "0" & shift_reg8 & shift_reg7 & shift_reg6 & shift_reg5 & shift_reg4 & shift_reg3 & shift_reg2 & shift_reg1);
	wire_add_sub5_datab <= ( "0" & shift_reg17 & shift_reg16 & shift_reg15 & shift_reg14 & shift_reg13 & shift_reg12 & shift_reg11 & shift_reg10);
	wire_add_sub5_w_result_range214w(0) <= wire_add_sub5_result(0);
	wire_add_sub5_w_result_range221w(0) <= wire_add_sub5_result(1);
	wire_add_sub5_w_result_range226w(0) <= wire_add_sub5_result(2);
	wire_add_sub5_w_result_range231w(0) <= wire_add_sub5_result(3);
	wire_add_sub5_w_result_range236w(0) <= wire_add_sub5_result(4);
	wire_add_sub5_w_result_range241w(0) <= wire_add_sub5_result(5);
	wire_add_sub5_w_result_range246w(0) <= wire_add_sub5_result(6);
	wire_add_sub5_w_result_range251w(0) <= wire_add_sub5_result(7);
	wire_add_sub5_w_result_range256w(0) <= wire_add_sub5_result(8);
	add_sub5 :  lpm_add_sub
	  GENERIC MAP (
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		cin => wire_gnd,
		dataa => wire_add_sub5_dataa,
		datab => wire_add_sub5_datab,
		result => wire_add_sub5_result
	  );
	wire_add_sub6_dataa <= ( data_in(8 DOWNTO 1));
	add_sub6 :  lpm_add_sub
	  GENERIC MAP (
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		cin => data_in(0),
		dataa => wire_add_sub6_dataa,
		result => wire_add_sub6_result
	  );
	wire_cmpr7_dataa <= ( data_in(7 DOWNTO 0));
	wire_cmpr7_datab <= "00000001";
	cmpr7 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aeb => wire_cmpr7_aeb,
		dataa => wire_cmpr7_dataa,
		datab => wire_cmpr7_datab
	  );
	cntr1 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "DOWN",
		lpm_modulus => 144,
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 8
	  )
	  PORT MAP ( 
		clock => clock,
		cnt_en => addr_counter_enable,
		data => addr_counter_sload_value,
		q => wire_cntr1_q,
		sload => addr_counter_sload
	  );
	cntr12 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "DOWN",
		lpm_modulus => 144,
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 8
	  )
	  PORT MAP ( 
		clock => clock,
		cnt_en => reconfig_addr_counter_enable,
		data => reconfig_addr_counter_sload_value,
		q => wire_cntr12_q,
		sload => reconfig_addr_counter_sload
	  );
	cntr13 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "DOWN",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 6
	  )
	  PORT MAP ( 
		clock => clock,
		cnt_en => reconfig_width_counter_enable,
		data => reconfig_width_counter_sload_value,
		q => wire_cntr13_q,
		sload => reconfig_width_counter_sload
	  );
	cntr14 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "DOWN",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 8
	  )
	  PORT MAP ( 
		clock => clock,
		cnt_en => rom_width_counter_enable,
		data => rom_width_counter_sload_value,
		q => wire_cntr14_q,
		sload => rom_width_counter_sload
	  );
	cntr15 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "DOWN",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 5
	  )
	  PORT MAP ( 
		clock => clock,
		cnt_en => rotate_width_counter_enable,
		data => rotate_width_counter_sload_value,
		q => wire_cntr15_q,
		sload => rotate_width_counter_sload
	  );
	cntr16 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "DOWN",
		lpm_modulus => 144,
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 8
	  )
	  PORT MAP ( 
		clock => clock,
		cnt_en => rotate_addr_counter_enable,
		data => rotate_addr_counter_sload_value,
		q => wire_cntr16_q,
		sload => rotate_addr_counter_sload
	  );
	cntr2 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 8
	  )
	  PORT MAP ( 
		clock => clock,
		cnt_en => read_addr_counter_enable,
		data => read_addr_counter_sload_value,
		q => wire_cntr2_q,
		sload => read_addr_counter_sload
	  );
	cntr3 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "DOWN",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 5
	  )
	  PORT MAP ( 
		clock => clock,
		cnt_en => width_counter_enable,
		data => width_counter_sload_value,
		q => wire_cntr3_q,
		sload => width_counter_sload
	  );
	decode11 :  lpm_decode
	  GENERIC MAP (
		LPM_DECODES => 5,
		LPM_WIDTH => 3
	  )
	  PORT MAP ( 
		data => cuda_combout_wire,
		eq => wire_decode11_eq
	  );

 END RTL; --video_pll_reconfig_pllrcfg_2871
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY video_pll_reconfig IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		counter_param		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		counter_type		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		data_in		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		pll_areset_in		: IN STD_LOGIC  := '0';
		pll_scandataout		: IN STD_LOGIC ;
		pll_scandone		: IN STD_LOGIC ;
		read_param		: IN STD_LOGIC ;
		reconfig		: IN STD_LOGIC ;
		reset		: IN STD_LOGIC ;
		reset_rom_address		: IN STD_LOGIC  := '0';
		rom_data_in		: IN STD_LOGIC  := '0';
		write_from_rom		: IN STD_LOGIC  := '0';
		write_param		: IN STD_LOGIC ;
		busy		: OUT STD_LOGIC ;
		data_out		: OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
		pll_areset		: OUT STD_LOGIC ;
		pll_configupdate		: OUT STD_LOGIC ;
		pll_scanclk		: OUT STD_LOGIC ;
		pll_scanclkena		: OUT STD_LOGIC ;
		pll_scandata		: OUT STD_LOGIC ;
		rom_address_out		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		write_rom_ena		: OUT STD_LOGIC 
	);
END video_pll_reconfig;


ARCHITECTURE RTL OF video_pll_reconfig IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "altpll_reconfig";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "init_from_external_rom_checkbox_checked=YES;init_from_rom=NO;intended_device_family=Cyclone 10 LP;scan_init_file=./Atari800XL/mist/ntsc.mif;";
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC ;
	SIGNAL sub_wire3	: STD_LOGIC ;
	SIGNAL sub_wire4	: STD_LOGIC ;
	SIGNAL sub_wire5	: STD_LOGIC ;
	SIGNAL sub_wire6	: STD_LOGIC ;
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC ;



	COMPONENT video_pll_reconfig_pllrcfg_2871
	PORT (
			clock	: IN STD_LOGIC ;
			counter_param	: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			counter_type	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			data_in	: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
			pll_areset_in	: IN STD_LOGIC ;
			pll_scandataout	: IN STD_LOGIC ;
			pll_scandone	: IN STD_LOGIC ;
			read_param	: IN STD_LOGIC ;
			reconfig	: IN STD_LOGIC ;
			reset	: IN STD_LOGIC ;
			reset_rom_address	: IN STD_LOGIC ;
			rom_data_in	: IN STD_LOGIC ;
			write_from_rom	: IN STD_LOGIC ;
			write_param	: IN STD_LOGIC ;
			busy	: OUT STD_LOGIC ;
			data_out	: OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
			pll_areset	: OUT STD_LOGIC ;
			pll_configupdate	: OUT STD_LOGIC ;
			pll_scanclk	: OUT STD_LOGIC ;
			pll_scanclkena	: OUT STD_LOGIC ;
			pll_scandata	: OUT STD_LOGIC ;
			rom_address_out	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			write_rom_ena	: OUT STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	busy    <= sub_wire0;
	data_out    <= sub_wire1(8 DOWNTO 0);
	pll_areset    <= sub_wire2;
	pll_configupdate    <= sub_wire3;
	pll_scanclk    <= sub_wire4;
	pll_scanclkena    <= sub_wire5;
	pll_scandata    <= sub_wire6;
	rom_address_out    <= sub_wire7(7 DOWNTO 0);
	write_rom_ena    <= sub_wire8;

	video_pll_reconfig_pllrcfg_2871_component : video_pll_reconfig_pllrcfg_2871
	PORT MAP (
		clock => clock,
		counter_param => counter_param,
		counter_type => counter_type,
		data_in => data_in,
		pll_areset_in => pll_areset_in,
		pll_scandataout => pll_scandataout,
		pll_scandone => pll_scandone,
		read_param => read_param,
		reconfig => reconfig,
		reset => reset,
		reset_rom_address => reset_rom_address,
		rom_data_in => rom_data_in,
		write_from_rom => write_from_rom,
		write_param => write_param,
		busy => sub_wire0,
		data_out => sub_wire1,
		pll_areset => sub_wire2,
		pll_configupdate => sub_wire3,
		pll_scanclk => sub_wire4,
		pll_scanclkena => sub_wire5,
		pll_scandata => sub_wire6,
		rom_address_out => sub_wire7,
		write_rom_ena => sub_wire8
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: CHAIN_TYPE NUMERIC "0"
-- Retrieval info: PRIVATE: INIT_FILE_NAME STRING "./Atari800XL/mist/ntsc.mif"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone 10 LP"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: USE_INIT_FILE STRING "1"
-- Retrieval info: CONSTANT: INIT_FROM_EXTERNAL_ROM_CHECKBOX_CHECKED STRING "YES"
-- Retrieval info: CONSTANT: INIT_FROM_ROM STRING "NO"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone 10 LP"
-- Retrieval info: CONSTANT: SCAN_INIT_FILE STRING "./Atari800XL/mist/ntsc.mif"
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: counter_param 0 0 3 0 INPUT NODEFVAL "counter_param[2..0]"
-- Retrieval info: USED_PORT: counter_type 0 0 4 0 INPUT NODEFVAL "counter_type[3..0]"
-- Retrieval info: USED_PORT: data_in 0 0 9 0 INPUT NODEFVAL "data_in[8..0]"
-- Retrieval info: USED_PORT: data_out 0 0 9 0 OUTPUT NODEFVAL "data_out[8..0]"
-- Retrieval info: USED_PORT: pll_areset 0 0 0 0 OUTPUT NODEFVAL "pll_areset"
-- Retrieval info: USED_PORT: pll_areset_in 0 0 0 0 INPUT GND "pll_areset_in"
-- Retrieval info: USED_PORT: pll_configupdate 0 0 0 0 OUTPUT NODEFVAL "pll_configupdate"
-- Retrieval info: USED_PORT: pll_scanclk 0 0 0 0 OUTPUT NODEFVAL "pll_scanclk"
-- Retrieval info: USED_PORT: pll_scanclkena 0 0 0 0 OUTPUT NODEFVAL "pll_scanclkena"
-- Retrieval info: USED_PORT: pll_scandata 0 0 0 0 OUTPUT NODEFVAL "pll_scandata"
-- Retrieval info: USED_PORT: pll_scandataout 0 0 0 0 INPUT NODEFVAL "pll_scandataout"
-- Retrieval info: USED_PORT: pll_scandone 0 0 0 0 INPUT NODEFVAL "pll_scandone"
-- Retrieval info: USED_PORT: read_param 0 0 0 0 INPUT NODEFVAL "read_param"
-- Retrieval info: USED_PORT: reconfig 0 0 0 0 INPUT NODEFVAL "reconfig"
-- Retrieval info: USED_PORT: reset 0 0 0 0 INPUT NODEFVAL "reset"
-- Retrieval info: USED_PORT: reset_rom_address 0 0 0 0 INPUT GND "reset_rom_address"
-- Retrieval info: USED_PORT: rom_address_out 0 0 8 0 OUTPUT NODEFVAL "rom_address_out[7..0]"
-- Retrieval info: USED_PORT: rom_data_in 0 0 0 0 INPUT GND "rom_data_in"
-- Retrieval info: USED_PORT: write_from_rom 0 0 0 0 INPUT GND "write_from_rom"
-- Retrieval info: USED_PORT: write_param 0 0 0 0 INPUT NODEFVAL "write_param"
-- Retrieval info: USED_PORT: write_rom_ena 0 0 0 0 OUTPUT NODEFVAL "write_rom_ena"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @counter_param 0 0 3 0 counter_param 0 0 3 0
-- Retrieval info: CONNECT: @counter_type 0 0 4 0 counter_type 0 0 4 0
-- Retrieval info: CONNECT: @data_in 0 0 9 0 data_in 0 0 9 0
-- Retrieval info: CONNECT: @pll_areset_in 0 0 0 0 pll_areset_in 0 0 0 0
-- Retrieval info: CONNECT: @pll_scandataout 0 0 0 0 pll_scandataout 0 0 0 0
-- Retrieval info: CONNECT: @pll_scandone 0 0 0 0 pll_scandone 0 0 0 0
-- Retrieval info: CONNECT: @read_param 0 0 0 0 read_param 0 0 0 0
-- Retrieval info: CONNECT: @reconfig 0 0 0 0 reconfig 0 0 0 0
-- Retrieval info: CONNECT: @reset 0 0 0 0 reset 0 0 0 0
-- Retrieval info: CONNECT: @reset_rom_address 0 0 0 0 reset_rom_address 0 0 0 0
-- Retrieval info: CONNECT: @rom_data_in 0 0 0 0 rom_data_in 0 0 0 0
-- Retrieval info: CONNECT: @write_from_rom 0 0 0 0 write_from_rom 0 0 0 0
-- Retrieval info: CONNECT: @write_param 0 0 0 0 write_param 0 0 0 0
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: CONNECT: data_out 0 0 9 0 @data_out 0 0 9 0
-- Retrieval info: CONNECT: pll_areset 0 0 0 0 @pll_areset 0 0 0 0
-- Retrieval info: CONNECT: pll_configupdate 0 0 0 0 @pll_configupdate 0 0 0 0
-- Retrieval info: CONNECT: pll_scanclk 0 0 0 0 @pll_scanclk 0 0 0 0
-- Retrieval info: CONNECT: pll_scanclkena 0 0 0 0 @pll_scanclkena 0 0 0 0
-- Retrieval info: CONNECT: pll_scandata 0 0 0 0 @pll_scandata 0 0 0 0
-- Retrieval info: CONNECT: rom_address_out 0 0 8 0 @rom_address_out 0 0 8 0
-- Retrieval info: CONNECT: write_rom_ena 0 0 0 0 @write_rom_ena 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL video_pll_reconfig.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL video_pll_reconfig.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL video_pll_reconfig.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL video_pll_reconfig.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL video_pll_reconfig_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
-- Retrieval info: LIB_FILE: cyclone10lp
-- Retrieval info: LIB_FILE: lpm
