
module pll_reconfig_calypso (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
